
module lpddr5_channel(
  clk,
  rst,
  read_clkEn,
  read_addr,
  read_req,
  read_busID,
  readOut_addr,
  readOut_req,
  readOut_busID,
  readOut_en,
  mem_clk,
  RAS,
  CAS,
  CS0,
  ADDR15,
  DATA18);
  parameter ODD_HALF=0;  
  
endmodule  
