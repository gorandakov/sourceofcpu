/*
Copyright 2022 Goran Dakov

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/


`include "../struct.sv"

module fprnd(
  A,
  rbit,tail,
  rndbit,
  rmode,
  isDBL,
  isEXT,
  toDBL,
  toSNG,
  B);
//rnd first, then denormal handling
  input [80:0] A;
  input rbit;
  input tail;
  input rndbit;
  input [2:0] rmode;
  input isDBL;
  input isEXT;
  input toDBL;
  input toSNG;
  output [79:0] B;

  wire [63:0] Ax;
  wire do_rnd;
  wire cout;

  assign Ax={A[63:53]&{11{isEXT}},A[52]|isDBL,A[51:0]};

  adder #(64) rnd_mod(Ax,rbit,res0,1'b0,do_rnd,cout);

  assign res0=~do_rnd ? Ax : 64'bz;
endmodule
