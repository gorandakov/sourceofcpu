
module insconv(
   bundle,
   bundle_out);

   input [255:0] bundle;
   output [255:0] bundle_out;

   wire [255:0] bundle_out_X; assign bundle_out=bundle_out_X;

   wire [14:-1] stp;

   assign bundle_out_X[239:0]=bundle[239:0];
   assign bundle_out_X[255]=bundle[255];

   assign stp={bundle[254:240],1'b1};

   generate
     genvar pos;
     for(pos=0;pos<15;pos=pos+1) begin
	 assign bundle_out_X[240+pos]=(stp[pos-1] && bundle[16*pos+:8]==8'hf2) || stp[pos];
     end
   endgenerate

endmodule
