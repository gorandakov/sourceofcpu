cntrl.cpp