
`define SR_FEXTCFG 64
`define SR_FDBLCFG 65


