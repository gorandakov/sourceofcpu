
`define mop_int8 3'd0
`define mop_int16 3'd1
`define mop_int32 3'd2
`define mop_int64 3'd3



