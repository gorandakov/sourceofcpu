  function [16:0] cnt0;
    input [15:0] bits;
    casex(bits)
        16'b0x0x0x0x0x0x0x0x : cnt0=17'h100;
        16'b10x0x0x0x0x0x0x0 : cnt0=17'h100;
        16'b110x0x0x0x0x0x0x : cnt0=17'h200;
        16'b0x10x0x0x0x0x0x0 : cnt0=17'h100;
        16'b1110x0x0x0x0x0x0 : cnt0=17'h200;
        16'b10x10x0x0x0x0x0x : cnt0=17'h200;
        16'b0x110x0x0x0x0x0x : cnt0=17'h200;
        16'b11110x0x0x0x0x0x : cnt0=17'h400;
        16'b0x0x10x0x0x0x0x0 : cnt0=17'h100;
        16'b110x10x0x0x0x0x0 : cnt0=17'h200;
        16'b10x110x0x0x0x0x0 : cnt0=17'h200;
        16'b0x1110x0x0x0x0x0 : cnt0=17'h200;
        16'b111110x0x0x0x0x0 : cnt0=17'h400;
        16'b10x0x10x0x0x0x0x : cnt0=17'h200;
        16'b0x10x10x0x0x0x0x : cnt0=17'h200;
        16'b1110x10x0x0x0x0x : cnt0=17'h400;
        16'b0x0x110x0x0x0x0x : cnt0=17'h200;
        16'b110x110x0x0x0x0x : cnt0=17'h400;
        16'b10x1110x0x0x0x0x : cnt0=17'h400;
        16'b0x11110x0x0x0x0x : cnt0=17'h400;
        16'b1111110x0x0x0x0x : cnt0=17'h800;
        16'b0x0x0x10x0x0x0x0 : cnt0=17'h100;
        16'b110x0x10x0x0x0x0 : cnt0=17'h200;
        16'b10x10x10x0x0x0x0 : cnt0=17'h200;
        16'b0x110x10x0x0x0x0 : cnt0=17'h200;
        16'b11110x10x0x0x0x0 : cnt0=17'h400;
        16'b10x0x110x0x0x0x0 : cnt0=17'h200;
        16'b0x10x110x0x0x0x0 : cnt0=17'h200;
        16'b1110x110x0x0x0x0 : cnt0=17'h400;
        16'b0x0x1110x0x0x0x0 : cnt0=17'h200;
        16'b110x1110x0x0x0x0 : cnt0=17'h400;
        16'b10x11110x0x0x0x0 : cnt0=17'h400;
        16'b0x111110x0x0x0x0 : cnt0=17'h400;
        16'b11111110x0x0x0x0 : cnt0=17'h800;
        16'b10x0x0x10x0x0x0x : cnt0=17'h200;
        16'b0x10x0x10x0x0x0x : cnt0=17'h200;
        16'b1110x0x10x0x0x0x : cnt0=17'h400;
        16'b0x0x10x10x0x0x0x : cnt0=17'h200;
        16'b110x10x10x0x0x0x : cnt0=17'h400;
        16'b10x110x10x0x0x0x : cnt0=17'h400;
        16'b0x1110x10x0x0x0x : cnt0=17'h400;
        16'b111110x10x0x0x0x : cnt0=17'h800;
        16'b0x0x0x110x0x0x0x : cnt0=17'h200;
        16'b110x0x110x0x0x0x : cnt0=17'h400;
        16'b10x10x110x0x0x0x : cnt0=17'h400;
        16'b0x110x110x0x0x0x : cnt0=17'h400;
        16'b11110x110x0x0x0x : cnt0=17'h800;
        16'b10x0x1110x0x0x0x : cnt0=17'h400;
        16'b0x10x1110x0x0x0x : cnt0=17'h400;
        16'b1110x1110x0x0x0x : cnt0=17'h800;
        16'b0x0x11110x0x0x0x : cnt0=17'h400;
        16'b110x11110x0x0x0x : cnt0=17'h800;
        16'b10x111110x0x0x0x : cnt0=17'h800;
        16'b0x1111110x0x0x0x : cnt0=17'h800;
        16'b111111110x0x0x0x : cnt0=17'h1000;
        16'b0x0x0x0x10x0x0x0 : cnt0=17'h100;
        16'b110x0x0x10x0x0x0 : cnt0=17'h200;
        16'b10x10x0x10x0x0x0 : cnt0=17'h200;
        16'b0x110x0x10x0x0x0 : cnt0=17'h200;
        16'b11110x0x10x0x0x0 : cnt0=17'h400;
        16'b10x0x10x10x0x0x0 : cnt0=17'h200;
        16'b0x10x10x10x0x0x0 : cnt0=17'h200;
        16'b1110x10x10x0x0x0 : cnt0=17'h400;
        16'b0x0x110x10x0x0x0 : cnt0=17'h200;
        16'b110x110x10x0x0x0 : cnt0=17'h400;
        16'b10x1110x10x0x0x0 : cnt0=17'h400;
        16'b0x11110x10x0x0x0 : cnt0=17'h400;
        16'b1111110x10x0x0x0 : cnt0=17'h800;
        16'b10x0x0x110x0x0x0 : cnt0=17'h200;
        16'b0x10x0x110x0x0x0 : cnt0=17'h200;
        16'b1110x0x110x0x0x0 : cnt0=17'h400;
        16'b0x0x10x110x0x0x0 : cnt0=17'h200;
        16'b110x10x110x0x0x0 : cnt0=17'h400;
        16'b10x110x110x0x0x0 : cnt0=17'h400;
        16'b0x1110x110x0x0x0 : cnt0=17'h400;
        16'b111110x110x0x0x0 : cnt0=17'h800;
        16'b0x0x0x1110x0x0x0 : cnt0=17'h200;
        16'b110x0x1110x0x0x0 : cnt0=17'h400;
        16'b10x10x1110x0x0x0 : cnt0=17'h400;
        16'b0x110x1110x0x0x0 : cnt0=17'h400;
        16'b11110x1110x0x0x0 : cnt0=17'h800;
        16'b10x0x11110x0x0x0 : cnt0=17'h400;
        16'b0x10x11110x0x0x0 : cnt0=17'h400;
        16'b1110x11110x0x0x0 : cnt0=17'h800;
        16'b0x0x111110x0x0x0 : cnt0=17'h400;
        16'b110x111110x0x0x0 : cnt0=17'h800;
        16'b10x1111110x0x0x0 : cnt0=17'h800;
        16'b0x11111110x0x0x0 : cnt0=17'h800;
        16'b1111111110x0x0x0 : cnt0=17'h1000;
        16'b10x0x0x0x10x0x0x : cnt0=17'h200;
        16'b0x10x0x0x10x0x0x : cnt0=17'h200;
        16'b1110x0x0x10x0x0x : cnt0=17'h400;
        16'b0x0x10x0x10x0x0x : cnt0=17'h200;
        16'b110x10x0x10x0x0x : cnt0=17'h400;
        16'b10x110x0x10x0x0x : cnt0=17'h400;
        16'b0x1110x0x10x0x0x : cnt0=17'h400;
        16'b111110x0x10x0x0x : cnt0=17'h800;
        16'b0x0x0x10x10x0x0x : cnt0=17'h200;
        16'b110x0x10x10x0x0x : cnt0=17'h400;
        16'b10x10x10x10x0x0x : cnt0=17'h400;
        16'b0x110x10x10x0x0x : cnt0=17'h400;
        16'b11110x10x10x0x0x : cnt0=17'h800;
        16'b10x0x110x10x0x0x : cnt0=17'h400;
        16'b0x10x110x10x0x0x : cnt0=17'h400;
        16'b1110x110x10x0x0x : cnt0=17'h800;
        16'b0x0x1110x10x0x0x : cnt0=17'h400;
        16'b110x1110x10x0x0x : cnt0=17'h800;
        16'b10x11110x10x0x0x : cnt0=17'h800;
        16'b0x111110x10x0x0x : cnt0=17'h800;
        16'b11111110x10x0x0x : cnt0=17'h1000;
        16'b0x0x0x0x110x0x0x : cnt0=17'h200;
        16'b110x0x0x110x0x0x : cnt0=17'h400;
        16'b10x10x0x110x0x0x : cnt0=17'h400;
        16'b0x110x0x110x0x0x : cnt0=17'h400;
        16'b11110x0x110x0x0x : cnt0=17'h800;
        16'b10x0x10x110x0x0x : cnt0=17'h400;
        16'b0x10x10x110x0x0x : cnt0=17'h400;
        16'b1110x10x110x0x0x : cnt0=17'h800;
        16'b0x0x110x110x0x0x : cnt0=17'h400;
        16'b110x110x110x0x0x : cnt0=17'h800;
        16'b10x1110x110x0x0x : cnt0=17'h800;
        16'b0x11110x110x0x0x : cnt0=17'h800;
        16'b1111110x110x0x0x : cnt0=17'h1000;
        16'b10x0x0x1110x0x0x : cnt0=17'h400;
        16'b0x10x0x1110x0x0x : cnt0=17'h400;
        16'b1110x0x1110x0x0x : cnt0=17'h800;
        16'b0x0x10x1110x0x0x : cnt0=17'h400;
        16'b110x10x1110x0x0x : cnt0=17'h800;
        16'b10x110x1110x0x0x : cnt0=17'h800;
        16'b0x1110x1110x0x0x : cnt0=17'h800;
        16'b111110x1110x0x0x : cnt0=17'h1000;
        16'b0x0x0x11110x0x0x : cnt0=17'h400;
        16'b110x0x11110x0x0x : cnt0=17'h800;
        16'b10x10x11110x0x0x : cnt0=17'h800;
        16'b0x110x11110x0x0x : cnt0=17'h800;
        16'b11110x11110x0x0x : cnt0=17'h1000;
        16'b10x0x111110x0x0x : cnt0=17'h800;
        16'b0x10x111110x0x0x : cnt0=17'h800;
        16'b1110x111110x0x0x : cnt0=17'h1000;
        16'b0x0x1111110x0x0x : cnt0=17'h800;
        16'b110x1111110x0x0x : cnt0=17'h1000;
        16'b10x11111110x0x0x : cnt0=17'h1000;
        16'b0x111111110x0x0x : cnt0=17'h1000;
        16'b11111111110x0x0x : cnt0=17'h2000;
        16'b0x0x0x0x0x10x0x0 : cnt0=17'h100;
        16'b110x0x0x0x10x0x0 : cnt0=17'h200;
        16'b10x10x0x0x10x0x0 : cnt0=17'h200;
        16'b0x110x0x0x10x0x0 : cnt0=17'h200;
        16'b11110x0x0x10x0x0 : cnt0=17'h400;
        16'b10x0x10x0x10x0x0 : cnt0=17'h200;
        16'b0x10x10x0x10x0x0 : cnt0=17'h200;
        16'b1110x10x0x10x0x0 : cnt0=17'h400;
        16'b0x0x110x0x10x0x0 : cnt0=17'h200;
        16'b110x110x0x10x0x0 : cnt0=17'h400;
        16'b10x1110x0x10x0x0 : cnt0=17'h400;
        16'b0x11110x0x10x0x0 : cnt0=17'h400;
        16'b1111110x0x10x0x0 : cnt0=17'h800;
        16'b10x0x0x10x10x0x0 : cnt0=17'h200;
        16'b0x10x0x10x10x0x0 : cnt0=17'h200;
        16'b1110x0x10x10x0x0 : cnt0=17'h400;
        16'b0x0x10x10x10x0x0 : cnt0=17'h200;
        16'b110x10x10x10x0x0 : cnt0=17'h400;
        16'b10x110x10x10x0x0 : cnt0=17'h400;
        16'b0x1110x10x10x0x0 : cnt0=17'h400;
        16'b111110x10x10x0x0 : cnt0=17'h800;
        16'b0x0x0x110x10x0x0 : cnt0=17'h200;
        16'b110x0x110x10x0x0 : cnt0=17'h400;
        16'b10x10x110x10x0x0 : cnt0=17'h400;
        16'b0x110x110x10x0x0 : cnt0=17'h400;
        16'b11110x110x10x0x0 : cnt0=17'h800;
        16'b10x0x1110x10x0x0 : cnt0=17'h400;
        16'b0x10x1110x10x0x0 : cnt0=17'h400;
        16'b1110x1110x10x0x0 : cnt0=17'h800;
        16'b0x0x11110x10x0x0 : cnt0=17'h400;
        16'b110x11110x10x0x0 : cnt0=17'h800;
        16'b10x111110x10x0x0 : cnt0=17'h800;
        16'b0x1111110x10x0x0 : cnt0=17'h800;
        16'b111111110x10x0x0 : cnt0=17'h1000;
        16'b10x0x0x0x110x0x0 : cnt0=17'h200;
        16'b0x10x0x0x110x0x0 : cnt0=17'h200;
        16'b1110x0x0x110x0x0 : cnt0=17'h400;
        16'b0x0x10x0x110x0x0 : cnt0=17'h200;
        16'b110x10x0x110x0x0 : cnt0=17'h400;
        16'b10x110x0x110x0x0 : cnt0=17'h400;
        16'b0x1110x0x110x0x0 : cnt0=17'h400;
        16'b111110x0x110x0x0 : cnt0=17'h800;
        16'b0x0x0x10x110x0x0 : cnt0=17'h200;
        16'b110x0x10x110x0x0 : cnt0=17'h400;
        16'b10x10x10x110x0x0 : cnt0=17'h400;
        16'b0x110x10x110x0x0 : cnt0=17'h400;
        16'b11110x10x110x0x0 : cnt0=17'h800;
        16'b10x0x110x110x0x0 : cnt0=17'h400;
        16'b0x10x110x110x0x0 : cnt0=17'h400;
        16'b1110x110x110x0x0 : cnt0=17'h800;
        16'b0x0x1110x110x0x0 : cnt0=17'h400;
        16'b110x1110x110x0x0 : cnt0=17'h800;
        16'b10x11110x110x0x0 : cnt0=17'h800;
        16'b0x111110x110x0x0 : cnt0=17'h800;
        16'b11111110x110x0x0 : cnt0=17'h1000;
        16'b0x0x0x0x1110x0x0 : cnt0=17'h200;
        16'b110x0x0x1110x0x0 : cnt0=17'h400;
        16'b10x10x0x1110x0x0 : cnt0=17'h400;
        16'b0x110x0x1110x0x0 : cnt0=17'h400;
        16'b11110x0x1110x0x0 : cnt0=17'h800;
        16'b10x0x10x1110x0x0 : cnt0=17'h400;
        16'b0x10x10x1110x0x0 : cnt0=17'h400;
        16'b1110x10x1110x0x0 : cnt0=17'h800;
        16'b0x0x110x1110x0x0 : cnt0=17'h400;
        16'b110x110x1110x0x0 : cnt0=17'h800;
        16'b10x1110x1110x0x0 : cnt0=17'h800;
        16'b0x11110x1110x0x0 : cnt0=17'h800;
        16'b1111110x1110x0x0 : cnt0=17'h1000;
        16'b10x0x0x11110x0x0 : cnt0=17'h400;
        16'b0x10x0x11110x0x0 : cnt0=17'h400;
        16'b1110x0x11110x0x0 : cnt0=17'h800;
        16'b0x0x10x11110x0x0 : cnt0=17'h400;
        16'b110x10x11110x0x0 : cnt0=17'h800;
        16'b10x110x11110x0x0 : cnt0=17'h800;
        16'b0x1110x11110x0x0 : cnt0=17'h800;
        16'b111110x11110x0x0 : cnt0=17'h1000;
        16'b0x0x0x111110x0x0 : cnt0=17'h400;
        16'b110x0x111110x0x0 : cnt0=17'h800;
        16'b10x10x111110x0x0 : cnt0=17'h800;
        16'b0x110x111110x0x0 : cnt0=17'h800;
        16'b11110x111110x0x0 : cnt0=17'h1000;
        16'b10x0x1111110x0x0 : cnt0=17'h800;
        16'b0x10x1111110x0x0 : cnt0=17'h800;
        16'b1110x1111110x0x0 : cnt0=17'h1000;
        16'b0x0x11111110x0x0 : cnt0=17'h800;
        16'b110x11111110x0x0 : cnt0=17'h1000;
        16'b10x111111110x0x0 : cnt0=17'h1000;
        16'b0x1111111110x0x0 : cnt0=17'h1000;
        16'b111111111110x0x0 : cnt0=17'h2000;
        16'b10x0x0x0x0x10x0x : cnt0=17'h200;
        16'b0x10x0x0x0x10x0x : cnt0=17'h200;
        16'b1110x0x0x0x10x0x : cnt0=17'h400;
        16'b0x0x10x0x0x10x0x : cnt0=17'h200;
        16'b110x10x0x0x10x0x : cnt0=17'h400;
        16'b10x110x0x0x10x0x : cnt0=17'h400;
        16'b0x1110x0x0x10x0x : cnt0=17'h400;
        16'b111110x0x0x10x0x : cnt0=17'h800;
        16'b0x0x0x10x0x10x0x : cnt0=17'h200;
        16'b110x0x10x0x10x0x : cnt0=17'h400;
        16'b10x10x10x0x10x0x : cnt0=17'h400;
        16'b0x110x10x0x10x0x : cnt0=17'h400;
        16'b11110x10x0x10x0x : cnt0=17'h800;
        16'b10x0x110x0x10x0x : cnt0=17'h400;
        16'b0x10x110x0x10x0x : cnt0=17'h400;
        16'b1110x110x0x10x0x : cnt0=17'h800;
        16'b0x0x1110x0x10x0x : cnt0=17'h400;
        16'b110x1110x0x10x0x : cnt0=17'h800;
        16'b10x11110x0x10x0x : cnt0=17'h800;
        16'b0x111110x0x10x0x : cnt0=17'h800;
        16'b11111110x0x10x0x : cnt0=17'h1000;
        16'b0x0x0x0x10x10x0x : cnt0=17'h200;
        16'b110x0x0x10x10x0x : cnt0=17'h400;
        16'b10x10x0x10x10x0x : cnt0=17'h400;
        16'b0x110x0x10x10x0x : cnt0=17'h400;
        16'b11110x0x10x10x0x : cnt0=17'h800;
        16'b10x0x10x10x10x0x : cnt0=17'h400;
        16'b0x10x10x10x10x0x : cnt0=17'h400;
        16'b1110x10x10x10x0x : cnt0=17'h800;
        16'b0x0x110x10x10x0x : cnt0=17'h400;
        16'b110x110x10x10x0x : cnt0=17'h800;
        16'b10x1110x10x10x0x : cnt0=17'h800;
        16'b0x11110x10x10x0x : cnt0=17'h800;
        16'b1111110x10x10x0x : cnt0=17'h1000;
        16'b10x0x0x110x10x0x : cnt0=17'h400;
        16'b0x10x0x110x10x0x : cnt0=17'h400;
        16'b1110x0x110x10x0x : cnt0=17'h800;
        16'b0x0x10x110x10x0x : cnt0=17'h400;
        16'b110x10x110x10x0x : cnt0=17'h800;
        16'b10x110x110x10x0x : cnt0=17'h800;
        16'b0x1110x110x10x0x : cnt0=17'h800;
        16'b111110x110x10x0x : cnt0=17'h1000;
        16'b0x0x0x1110x10x0x : cnt0=17'h400;
        16'b110x0x1110x10x0x : cnt0=17'h800;
        16'b10x10x1110x10x0x : cnt0=17'h800;
        16'b0x110x1110x10x0x : cnt0=17'h800;
        16'b11110x1110x10x0x : cnt0=17'h1000;
        16'b10x0x11110x10x0x : cnt0=17'h800;
        16'b0x10x11110x10x0x : cnt0=17'h800;
        16'b1110x11110x10x0x : cnt0=17'h1000;
        16'b0x0x111110x10x0x : cnt0=17'h800;
        16'b110x111110x10x0x : cnt0=17'h1000;
        16'b10x1111110x10x0x : cnt0=17'h1000;
        16'b0x11111110x10x0x : cnt0=17'h1000;
        16'b1111111110x10x0x : cnt0=17'h2000;
        16'b0x0x0x0x0x110x0x : cnt0=17'h200;
        16'b110x0x0x0x110x0x : cnt0=17'h400;
        16'b10x10x0x0x110x0x : cnt0=17'h400;
        16'b0x110x0x0x110x0x : cnt0=17'h400;
        16'b11110x0x0x110x0x : cnt0=17'h800;
        16'b10x0x10x0x110x0x : cnt0=17'h400;
        16'b0x10x10x0x110x0x : cnt0=17'h400;
        16'b1110x10x0x110x0x : cnt0=17'h800;
        16'b0x0x110x0x110x0x : cnt0=17'h400;
        16'b110x110x0x110x0x : cnt0=17'h800;
        16'b10x1110x0x110x0x : cnt0=17'h800;
        16'b0x11110x0x110x0x : cnt0=17'h800;
        16'b1111110x0x110x0x : cnt0=17'h1000;
        16'b10x0x0x10x110x0x : cnt0=17'h400;
        16'b0x10x0x10x110x0x : cnt0=17'h400;
        16'b1110x0x10x110x0x : cnt0=17'h800;
        16'b0x0x10x10x110x0x : cnt0=17'h400;
        16'b110x10x10x110x0x : cnt0=17'h800;
        16'b10x110x10x110x0x : cnt0=17'h800;
        16'b0x1110x10x110x0x : cnt0=17'h800;
        16'b111110x10x110x0x : cnt0=17'h1000;
        16'b0x0x0x110x110x0x : cnt0=17'h400;
        16'b110x0x110x110x0x : cnt0=17'h800;
        16'b10x10x110x110x0x : cnt0=17'h800;
        16'b0x110x110x110x0x : cnt0=17'h800;
        16'b11110x110x110x0x : cnt0=17'h1000;
        16'b10x0x1110x110x0x : cnt0=17'h800;
        16'b0x10x1110x110x0x : cnt0=17'h800;
        16'b1110x1110x110x0x : cnt0=17'h1000;
        16'b0x0x11110x110x0x : cnt0=17'h800;
        16'b110x11110x110x0x : cnt0=17'h1000;
        16'b10x111110x110x0x : cnt0=17'h1000;
        16'b0x1111110x110x0x : cnt0=17'h1000;
        16'b111111110x110x0x : cnt0=17'h2000;
        16'b10x0x0x0x1110x0x : cnt0=17'h400;
        16'b0x10x0x0x1110x0x : cnt0=17'h400;
        16'b1110x0x0x1110x0x : cnt0=17'h800;
        16'b0x0x10x0x1110x0x : cnt0=17'h400;
        16'b110x10x0x1110x0x : cnt0=17'h800;
        16'b10x110x0x1110x0x : cnt0=17'h800;
        16'b0x1110x0x1110x0x : cnt0=17'h800;
        16'b111110x0x1110x0x : cnt0=17'h1000;
        16'b0x0x0x10x1110x0x : cnt0=17'h400;
        16'b110x0x10x1110x0x : cnt0=17'h800;
        16'b10x10x10x1110x0x : cnt0=17'h800;
        16'b0x110x10x1110x0x : cnt0=17'h800;
        16'b11110x10x1110x0x : cnt0=17'h1000;
        16'b10x0x110x1110x0x : cnt0=17'h800;
        16'b0x10x110x1110x0x : cnt0=17'h800;
        16'b1110x110x1110x0x : cnt0=17'h1000;
        16'b0x0x1110x1110x0x : cnt0=17'h800;
        16'b110x1110x1110x0x : cnt0=17'h1000;
        16'b10x11110x1110x0x : cnt0=17'h1000;
        16'b0x111110x1110x0x : cnt0=17'h1000;
        16'b11111110x1110x0x : cnt0=17'h2000;
        16'b0x0x0x0x11110x0x : cnt0=17'h400;
        16'b110x0x0x11110x0x : cnt0=17'h800;
        16'b10x10x0x11110x0x : cnt0=17'h800;
        16'b0x110x0x11110x0x : cnt0=17'h800;
        16'b11110x0x11110x0x : cnt0=17'h1000;
        16'b10x0x10x11110x0x : cnt0=17'h800;
        16'b0x10x10x11110x0x : cnt0=17'h800;
        16'b1110x10x11110x0x : cnt0=17'h1000;
        16'b0x0x110x11110x0x : cnt0=17'h800;
        16'b110x110x11110x0x : cnt0=17'h1000;
        16'b10x1110x11110x0x : cnt0=17'h1000;
        16'b0x11110x11110x0x : cnt0=17'h1000;
        16'b1111110x11110x0x : cnt0=17'h2000;
        16'b10x0x0x111110x0x : cnt0=17'h800;
        16'b0x10x0x111110x0x : cnt0=17'h800;
        16'b1110x0x111110x0x : cnt0=17'h1000;
        16'b0x0x10x111110x0x : cnt0=17'h800;
        16'b110x10x111110x0x : cnt0=17'h1000;
        16'b10x110x111110x0x : cnt0=17'h1000;
        16'b0x1110x111110x0x : cnt0=17'h1000;
        16'b111110x111110x0x : cnt0=17'h2000;
        16'b0x0x0x1111110x0x : cnt0=17'h800;
        16'b110x0x1111110x0x : cnt0=17'h1000;
        16'b10x10x1111110x0x : cnt0=17'h1000;
        16'b0x110x1111110x0x : cnt0=17'h1000;
        16'b11110x1111110x0x : cnt0=17'h2000;
        16'b10x0x11111110x0x : cnt0=17'h1000;
        16'b0x10x11111110x0x : cnt0=17'h1000;
        16'b1110x11111110x0x : cnt0=17'h2000;
        16'b0x0x111111110x0x : cnt0=17'h1000;
        16'b110x111111110x0x : cnt0=17'h2000;
        16'b10x1111111110x0x : cnt0=17'h2000;
        16'b0x11111111110x0x : cnt0=17'h2000;
        16'b1111111111110x0x : cnt0=17'h4000;
        16'b0x0x0x0x0x0x10x0 : cnt0=17'h100;
        16'b110x0x0x0x0x10x0 : cnt0=17'h200;
        16'b10x10x0x0x0x10x0 : cnt0=17'h200;
        16'b0x110x0x0x0x10x0 : cnt0=17'h200;
        16'b11110x0x0x0x10x0 : cnt0=17'h400;
        16'b10x0x10x0x0x10x0 : cnt0=17'h200;
        16'b0x10x10x0x0x10x0 : cnt0=17'h200;
        16'b1110x10x0x0x10x0 : cnt0=17'h400;
        16'b0x0x110x0x0x10x0 : cnt0=17'h200;
        16'b110x110x0x0x10x0 : cnt0=17'h400;
        16'b10x1110x0x0x10x0 : cnt0=17'h400;
        16'b0x11110x0x0x10x0 : cnt0=17'h400;
        16'b1111110x0x0x10x0 : cnt0=17'h800;
        16'b10x0x0x10x0x10x0 : cnt0=17'h200;
        16'b0x10x0x10x0x10x0 : cnt0=17'h200;
        16'b1110x0x10x0x10x0 : cnt0=17'h400;
        16'b0x0x10x10x0x10x0 : cnt0=17'h200;
        16'b110x10x10x0x10x0 : cnt0=17'h400;
        16'b10x110x10x0x10x0 : cnt0=17'h400;
        16'b0x1110x10x0x10x0 : cnt0=17'h400;
        16'b111110x10x0x10x0 : cnt0=17'h800;
        16'b0x0x0x110x0x10x0 : cnt0=17'h200;
        16'b110x0x110x0x10x0 : cnt0=17'h400;
        16'b10x10x110x0x10x0 : cnt0=17'h400;
        16'b0x110x110x0x10x0 : cnt0=17'h400;
        16'b11110x110x0x10x0 : cnt0=17'h800;
        16'b10x0x1110x0x10x0 : cnt0=17'h400;
        16'b0x10x1110x0x10x0 : cnt0=17'h400;
        16'b1110x1110x0x10x0 : cnt0=17'h800;
        16'b0x0x11110x0x10x0 : cnt0=17'h400;
        16'b110x11110x0x10x0 : cnt0=17'h800;
        16'b10x111110x0x10x0 : cnt0=17'h800;
        16'b0x1111110x0x10x0 : cnt0=17'h800;
        16'b111111110x0x10x0 : cnt0=17'h1000;
        16'b10x0x0x0x10x10x0 : cnt0=17'h200;
        16'b0x10x0x0x10x10x0 : cnt0=17'h200;
        16'b1110x0x0x10x10x0 : cnt0=17'h400;
        16'b0x0x10x0x10x10x0 : cnt0=17'h200;
        16'b110x10x0x10x10x0 : cnt0=17'h400;
        16'b10x110x0x10x10x0 : cnt0=17'h400;
        16'b0x1110x0x10x10x0 : cnt0=17'h400;
        16'b111110x0x10x10x0 : cnt0=17'h800;
        16'b0x0x0x10x10x10x0 : cnt0=17'h200;
        16'b110x0x10x10x10x0 : cnt0=17'h400;
        16'b10x10x10x10x10x0 : cnt0=17'h400;
        16'b0x110x10x10x10x0 : cnt0=17'h400;
        16'b11110x10x10x10x0 : cnt0=17'h800;
        16'b10x0x110x10x10x0 : cnt0=17'h400;
        16'b0x10x110x10x10x0 : cnt0=17'h400;
        16'b1110x110x10x10x0 : cnt0=17'h800;
        16'b0x0x1110x10x10x0 : cnt0=17'h400;
        16'b110x1110x10x10x0 : cnt0=17'h800;
        16'b10x11110x10x10x0 : cnt0=17'h800;
        16'b0x111110x10x10x0 : cnt0=17'h800;
        16'b11111110x10x10x0 : cnt0=17'h1000;
        16'b0x0x0x0x110x10x0 : cnt0=17'h200;
        16'b110x0x0x110x10x0 : cnt0=17'h400;
        16'b10x10x0x110x10x0 : cnt0=17'h400;
        16'b0x110x0x110x10x0 : cnt0=17'h400;
        16'b11110x0x110x10x0 : cnt0=17'h800;
        16'b10x0x10x110x10x0 : cnt0=17'h400;
        16'b0x10x10x110x10x0 : cnt0=17'h400;
        16'b1110x10x110x10x0 : cnt0=17'h800;
        16'b0x0x110x110x10x0 : cnt0=17'h400;
        16'b110x110x110x10x0 : cnt0=17'h800;
        16'b10x1110x110x10x0 : cnt0=17'h800;
        16'b0x11110x110x10x0 : cnt0=17'h800;
        16'b1111110x110x10x0 : cnt0=17'h1000;
        16'b10x0x0x1110x10x0 : cnt0=17'h400;
        16'b0x10x0x1110x10x0 : cnt0=17'h400;
        16'b1110x0x1110x10x0 : cnt0=17'h800;
        16'b0x0x10x1110x10x0 : cnt0=17'h400;
        16'b110x10x1110x10x0 : cnt0=17'h800;
        16'b10x110x1110x10x0 : cnt0=17'h800;
        16'b0x1110x1110x10x0 : cnt0=17'h800;
        16'b111110x1110x10x0 : cnt0=17'h1000;
        16'b0x0x0x11110x10x0 : cnt0=17'h400;
        16'b110x0x11110x10x0 : cnt0=17'h800;
        16'b10x10x11110x10x0 : cnt0=17'h800;
        16'b0x110x11110x10x0 : cnt0=17'h800;
        16'b11110x11110x10x0 : cnt0=17'h1000;
        16'b10x0x111110x10x0 : cnt0=17'h800;
        16'b0x10x111110x10x0 : cnt0=17'h800;
        16'b1110x111110x10x0 : cnt0=17'h1000;
        16'b0x0x1111110x10x0 : cnt0=17'h800;
        16'b110x1111110x10x0 : cnt0=17'h1000;
        16'b10x11111110x10x0 : cnt0=17'h1000;
        16'b0x111111110x10x0 : cnt0=17'h1000;
        16'b11111111110x10x0 : cnt0=17'h2000;
        16'b10x0x0x0x0x110x0 : cnt0=17'h200;
        16'b0x10x0x0x0x110x0 : cnt0=17'h200;
        16'b1110x0x0x0x110x0 : cnt0=17'h400;
        16'b0x0x10x0x0x110x0 : cnt0=17'h200;
        16'b110x10x0x0x110x0 : cnt0=17'h400;
        16'b10x110x0x0x110x0 : cnt0=17'h400;
        16'b0x1110x0x0x110x0 : cnt0=17'h400;
        16'b111110x0x0x110x0 : cnt0=17'h800;
        16'b0x0x0x10x0x110x0 : cnt0=17'h200;
        16'b110x0x10x0x110x0 : cnt0=17'h400;
        16'b10x10x10x0x110x0 : cnt0=17'h400;
        16'b0x110x10x0x110x0 : cnt0=17'h400;
        16'b11110x10x0x110x0 : cnt0=17'h800;
        16'b10x0x110x0x110x0 : cnt0=17'h400;
        16'b0x10x110x0x110x0 : cnt0=17'h400;
        16'b1110x110x0x110x0 : cnt0=17'h800;
        16'b0x0x1110x0x110x0 : cnt0=17'h400;
        16'b110x1110x0x110x0 : cnt0=17'h800;
        16'b10x11110x0x110x0 : cnt0=17'h800;
        16'b0x111110x0x110x0 : cnt0=17'h800;
        16'b11111110x0x110x0 : cnt0=17'h1000;
        16'b0x0x0x0x10x110x0 : cnt0=17'h200;
        16'b110x0x0x10x110x0 : cnt0=17'h400;
        16'b10x10x0x10x110x0 : cnt0=17'h400;
        16'b0x110x0x10x110x0 : cnt0=17'h400;
        16'b11110x0x10x110x0 : cnt0=17'h800;
        16'b10x0x10x10x110x0 : cnt0=17'h400;
        16'b0x10x10x10x110x0 : cnt0=17'h400;
        16'b1110x10x10x110x0 : cnt0=17'h800;
        16'b0x0x110x10x110x0 : cnt0=17'h400;
        16'b110x110x10x110x0 : cnt0=17'h800;
        16'b10x1110x10x110x0 : cnt0=17'h800;
        16'b0x11110x10x110x0 : cnt0=17'h800;
        16'b1111110x10x110x0 : cnt0=17'h1000;
        16'b10x0x0x110x110x0 : cnt0=17'h400;
        16'b0x10x0x110x110x0 : cnt0=17'h400;
        16'b1110x0x110x110x0 : cnt0=17'h800;
        16'b0x0x10x110x110x0 : cnt0=17'h400;
        16'b110x10x110x110x0 : cnt0=17'h800;
        16'b10x110x110x110x0 : cnt0=17'h800;
        16'b0x1110x110x110x0 : cnt0=17'h800;
        16'b111110x110x110x0 : cnt0=17'h1000;
        16'b0x0x0x1110x110x0 : cnt0=17'h400;
        16'b110x0x1110x110x0 : cnt0=17'h800;
        16'b10x10x1110x110x0 : cnt0=17'h800;
        16'b0x110x1110x110x0 : cnt0=17'h800;
        16'b11110x1110x110x0 : cnt0=17'h1000;
        16'b10x0x11110x110x0 : cnt0=17'h800;
        16'b0x10x11110x110x0 : cnt0=17'h800;
        16'b1110x11110x110x0 : cnt0=17'h1000;
        16'b0x0x111110x110x0 : cnt0=17'h800;
        16'b110x111110x110x0 : cnt0=17'h1000;
        16'b10x1111110x110x0 : cnt0=17'h1000;
        16'b0x11111110x110x0 : cnt0=17'h1000;
        16'b1111111110x110x0 : cnt0=17'h2000;
        16'b0x0x0x0x0x1110x0 : cnt0=17'h200;
        16'b110x0x0x0x1110x0 : cnt0=17'h400;
        16'b10x10x0x0x1110x0 : cnt0=17'h400;
        16'b0x110x0x0x1110x0 : cnt0=17'h400;
        16'b11110x0x0x1110x0 : cnt0=17'h800;
        16'b10x0x10x0x1110x0 : cnt0=17'h400;
        16'b0x10x10x0x1110x0 : cnt0=17'h400;
        16'b1110x10x0x1110x0 : cnt0=17'h800;
        16'b0x0x110x0x1110x0 : cnt0=17'h400;
        16'b110x110x0x1110x0 : cnt0=17'h800;
        16'b10x1110x0x1110x0 : cnt0=17'h800;
        16'b0x11110x0x1110x0 : cnt0=17'h800;
        16'b1111110x0x1110x0 : cnt0=17'h1000;
        16'b10x0x0x10x1110x0 : cnt0=17'h400;
        16'b0x10x0x10x1110x0 : cnt0=17'h400;
        16'b1110x0x10x1110x0 : cnt0=17'h800;
        16'b0x0x10x10x1110x0 : cnt0=17'h400;
        16'b110x10x10x1110x0 : cnt0=17'h800;
        16'b10x110x10x1110x0 : cnt0=17'h800;
        16'b0x1110x10x1110x0 : cnt0=17'h800;
        16'b111110x10x1110x0 : cnt0=17'h1000;
        16'b0x0x0x110x1110x0 : cnt0=17'h400;
        16'b110x0x110x1110x0 : cnt0=17'h800;
        16'b10x10x110x1110x0 : cnt0=17'h800;
        16'b0x110x110x1110x0 : cnt0=17'h800;
        16'b11110x110x1110x0 : cnt0=17'h1000;
        16'b10x0x1110x1110x0 : cnt0=17'h800;
        16'b0x10x1110x1110x0 : cnt0=17'h800;
        16'b1110x1110x1110x0 : cnt0=17'h1000;
        16'b0x0x11110x1110x0 : cnt0=17'h800;
        16'b110x11110x1110x0 : cnt0=17'h1000;
        16'b10x111110x1110x0 : cnt0=17'h1000;
        16'b0x1111110x1110x0 : cnt0=17'h1000;
        16'b111111110x1110x0 : cnt0=17'h2000;
        16'b10x0x0x0x11110x0 : cnt0=17'h400;
        16'b0x10x0x0x11110x0 : cnt0=17'h400;
        16'b1110x0x0x11110x0 : cnt0=17'h800;
        16'b0x0x10x0x11110x0 : cnt0=17'h400;
        16'b110x10x0x11110x0 : cnt0=17'h800;
        16'b10x110x0x11110x0 : cnt0=17'h800;
        16'b0x1110x0x11110x0 : cnt0=17'h800;
        16'b111110x0x11110x0 : cnt0=17'h1000;
        16'b0x0x0x10x11110x0 : cnt0=17'h400;
        16'b110x0x10x11110x0 : cnt0=17'h800;
        16'b10x10x10x11110x0 : cnt0=17'h800;
        16'b0x110x10x11110x0 : cnt0=17'h800;
        16'b11110x10x11110x0 : cnt0=17'h1000;
        16'b10x0x110x11110x0 : cnt0=17'h800;
        16'b0x10x110x11110x0 : cnt0=17'h800;
        16'b1110x110x11110x0 : cnt0=17'h1000;
        16'b0x0x1110x11110x0 : cnt0=17'h800;
        16'b110x1110x11110x0 : cnt0=17'h1000;
        16'b10x11110x11110x0 : cnt0=17'h1000;
        16'b0x111110x11110x0 : cnt0=17'h1000;
        16'b11111110x11110x0 : cnt0=17'h2000;
        16'b0x0x0x0x111110x0 : cnt0=17'h400;
        16'b110x0x0x111110x0 : cnt0=17'h800;
        16'b10x10x0x111110x0 : cnt0=17'h800;
        16'b0x110x0x111110x0 : cnt0=17'h800;
        16'b11110x0x111110x0 : cnt0=17'h1000;
        16'b10x0x10x111110x0 : cnt0=17'h800;
        16'b0x10x10x111110x0 : cnt0=17'h800;
        16'b1110x10x111110x0 : cnt0=17'h1000;
        16'b0x0x110x111110x0 : cnt0=17'h800;
        16'b110x110x111110x0 : cnt0=17'h1000;
        16'b10x1110x111110x0 : cnt0=17'h1000;
        16'b0x11110x111110x0 : cnt0=17'h1000;
        16'b1111110x111110x0 : cnt0=17'h2000;
        16'b10x0x0x1111110x0 : cnt0=17'h800;
        16'b0x10x0x1111110x0 : cnt0=17'h800;
        16'b1110x0x1111110x0 : cnt0=17'h1000;
        16'b0x0x10x1111110x0 : cnt0=17'h800;
        16'b110x10x1111110x0 : cnt0=17'h1000;
        16'b10x110x1111110x0 : cnt0=17'h1000;
        16'b0x1110x1111110x0 : cnt0=17'h1000;
        16'b111110x1111110x0 : cnt0=17'h2000;
        16'b0x0x0x11111110x0 : cnt0=17'h800;
        16'b110x0x11111110x0 : cnt0=17'h1000;
        16'b10x10x11111110x0 : cnt0=17'h1000;
        16'b0x110x11111110x0 : cnt0=17'h1000;
        16'b11110x11111110x0 : cnt0=17'h2000;
        16'b10x0x111111110x0 : cnt0=17'h1000;
        16'b0x10x111111110x0 : cnt0=17'h1000;
        16'b1110x111111110x0 : cnt0=17'h2000;
        16'b0x0x1111111110x0 : cnt0=17'h1000;
        16'b110x1111111110x0 : cnt0=17'h2000;
        16'b10x11111111110x0 : cnt0=17'h2000;
        16'b0x111111111110x0 : cnt0=17'h2000;
        16'b11111111111110x0 : cnt0=17'h4000;
        16'b10x0x0x0x0x0x10x : cnt0=17'h200;
        16'b0x10x0x0x0x0x10x : cnt0=17'h200;
        16'b1110x0x0x0x0x10x : cnt0=17'h400;
        16'b0x0x10x0x0x0x10x : cnt0=17'h200;
        16'b110x10x0x0x0x10x : cnt0=17'h400;
        16'b10x110x0x0x0x10x : cnt0=17'h400;
        16'b0x1110x0x0x0x10x : cnt0=17'h400;
        16'b111110x0x0x0x10x : cnt0=17'h800;
        16'b0x0x0x10x0x0x10x : cnt0=17'h200;
        16'b110x0x10x0x0x10x : cnt0=17'h400;
        16'b10x10x10x0x0x10x : cnt0=17'h400;
        16'b0x110x10x0x0x10x : cnt0=17'h400;
        16'b11110x10x0x0x10x : cnt0=17'h800;
        16'b10x0x110x0x0x10x : cnt0=17'h400;
        16'b0x10x110x0x0x10x : cnt0=17'h400;
        16'b1110x110x0x0x10x : cnt0=17'h800;
        16'b0x0x1110x0x0x10x : cnt0=17'h400;
        16'b110x1110x0x0x10x : cnt0=17'h800;
        16'b10x11110x0x0x10x : cnt0=17'h800;
        16'b0x111110x0x0x10x : cnt0=17'h800;
        16'b11111110x0x0x10x : cnt0=17'h1000;
        16'b0x0x0x0x10x0x10x : cnt0=17'h200;
        16'b110x0x0x10x0x10x : cnt0=17'h400;
        16'b10x10x0x10x0x10x : cnt0=17'h400;
        16'b0x110x0x10x0x10x : cnt0=17'h400;
        16'b11110x0x10x0x10x : cnt0=17'h800;
        16'b10x0x10x10x0x10x : cnt0=17'h400;
        16'b0x10x10x10x0x10x : cnt0=17'h400;
        16'b1110x10x10x0x10x : cnt0=17'h800;
        16'b0x0x110x10x0x10x : cnt0=17'h400;
        16'b110x110x10x0x10x : cnt0=17'h800;
        16'b10x1110x10x0x10x : cnt0=17'h800;
        16'b0x11110x10x0x10x : cnt0=17'h800;
        16'b1111110x10x0x10x : cnt0=17'h1000;
        16'b10x0x0x110x0x10x : cnt0=17'h400;
        16'b0x10x0x110x0x10x : cnt0=17'h400;
        16'b1110x0x110x0x10x : cnt0=17'h800;
        16'b0x0x10x110x0x10x : cnt0=17'h400;
        16'b110x10x110x0x10x : cnt0=17'h800;
        16'b10x110x110x0x10x : cnt0=17'h800;
        16'b0x1110x110x0x10x : cnt0=17'h800;
        16'b111110x110x0x10x : cnt0=17'h1000;
        16'b0x0x0x1110x0x10x : cnt0=17'h400;
        16'b110x0x1110x0x10x : cnt0=17'h800;
        16'b10x10x1110x0x10x : cnt0=17'h800;
        16'b0x110x1110x0x10x : cnt0=17'h800;
        16'b11110x1110x0x10x : cnt0=17'h1000;
        16'b10x0x11110x0x10x : cnt0=17'h800;
        16'b0x10x11110x0x10x : cnt0=17'h800;
        16'b1110x11110x0x10x : cnt0=17'h1000;
        16'b0x0x111110x0x10x : cnt0=17'h800;
        16'b110x111110x0x10x : cnt0=17'h1000;
        16'b10x1111110x0x10x : cnt0=17'h1000;
        16'b0x11111110x0x10x : cnt0=17'h1000;
        16'b1111111110x0x10x : cnt0=17'h2000;
        16'b0x0x0x0x0x10x10x : cnt0=17'h200;
        16'b110x0x0x0x10x10x : cnt0=17'h400;
        16'b10x10x0x0x10x10x : cnt0=17'h400;
        16'b0x110x0x0x10x10x : cnt0=17'h400;
        16'b11110x0x0x10x10x : cnt0=17'h800;
        16'b10x0x10x0x10x10x : cnt0=17'h400;
        16'b0x10x10x0x10x10x : cnt0=17'h400;
        16'b1110x10x0x10x10x : cnt0=17'h800;
        16'b0x0x110x0x10x10x : cnt0=17'h400;
        16'b110x110x0x10x10x : cnt0=17'h800;
        16'b10x1110x0x10x10x : cnt0=17'h800;
        16'b0x11110x0x10x10x : cnt0=17'h800;
        16'b1111110x0x10x10x : cnt0=17'h1000;
        16'b10x0x0x10x10x10x : cnt0=17'h400;
        16'b0x10x0x10x10x10x : cnt0=17'h400;
        16'b1110x0x10x10x10x : cnt0=17'h800;
        16'b0x0x10x10x10x10x : cnt0=17'h400;
        16'b110x10x10x10x10x : cnt0=17'h800;
        16'b10x110x10x10x10x : cnt0=17'h800;
        16'b0x1110x10x10x10x : cnt0=17'h800;
        16'b111110x10x10x10x : cnt0=17'h1000;
        16'b0x0x0x110x10x10x : cnt0=17'h400;
        16'b110x0x110x10x10x : cnt0=17'h800;
        16'b10x10x110x10x10x : cnt0=17'h800;
        16'b0x110x110x10x10x : cnt0=17'h800;
        16'b11110x110x10x10x : cnt0=17'h1000;
        16'b10x0x1110x10x10x : cnt0=17'h800;
        16'b0x10x1110x10x10x : cnt0=17'h800;
        16'b1110x1110x10x10x : cnt0=17'h1000;
        16'b0x0x11110x10x10x : cnt0=17'h800;
        16'b110x11110x10x10x : cnt0=17'h1000;
        16'b10x111110x10x10x : cnt0=17'h1000;
        16'b0x1111110x10x10x : cnt0=17'h1000;
        16'b111111110x10x10x : cnt0=17'h2000;
        16'b10x0x0x0x110x10x : cnt0=17'h400;
        16'b0x10x0x0x110x10x : cnt0=17'h400;
        16'b1110x0x0x110x10x : cnt0=17'h800;
        16'b0x0x10x0x110x10x : cnt0=17'h400;
        16'b110x10x0x110x10x : cnt0=17'h800;
        16'b10x110x0x110x10x : cnt0=17'h800;
        16'b0x1110x0x110x10x : cnt0=17'h800;
        16'b111110x0x110x10x : cnt0=17'h1000;
        16'b0x0x0x10x110x10x : cnt0=17'h400;
        16'b110x0x10x110x10x : cnt0=17'h800;
        16'b10x10x10x110x10x : cnt0=17'h800;
        16'b0x110x10x110x10x : cnt0=17'h800;
        16'b11110x10x110x10x : cnt0=17'h1000;
        16'b10x0x110x110x10x : cnt0=17'h800;
        16'b0x10x110x110x10x : cnt0=17'h800;
        16'b1110x110x110x10x : cnt0=17'h1000;
        16'b0x0x1110x110x10x : cnt0=17'h800;
        16'b110x1110x110x10x : cnt0=17'h1000;
        16'b10x11110x110x10x : cnt0=17'h1000;
        16'b0x111110x110x10x : cnt0=17'h1000;
        16'b11111110x110x10x : cnt0=17'h2000;
        16'b0x0x0x0x1110x10x : cnt0=17'h400;
        16'b110x0x0x1110x10x : cnt0=17'h800;
        16'b10x10x0x1110x10x : cnt0=17'h800;
        16'b0x110x0x1110x10x : cnt0=17'h800;
        16'b11110x0x1110x10x : cnt0=17'h1000;
        16'b10x0x10x1110x10x : cnt0=17'h800;
        16'b0x10x10x1110x10x : cnt0=17'h800;
        16'b1110x10x1110x10x : cnt0=17'h1000;
        16'b0x0x110x1110x10x : cnt0=17'h800;
        16'b110x110x1110x10x : cnt0=17'h1000;
        16'b10x1110x1110x10x : cnt0=17'h1000;
        16'b0x11110x1110x10x : cnt0=17'h1000;
        16'b1111110x1110x10x : cnt0=17'h2000;
        16'b10x0x0x11110x10x : cnt0=17'h800;
        16'b0x10x0x11110x10x : cnt0=17'h800;
        16'b1110x0x11110x10x : cnt0=17'h1000;
        16'b0x0x10x11110x10x : cnt0=17'h800;
        16'b110x10x11110x10x : cnt0=17'h1000;
        16'b10x110x11110x10x : cnt0=17'h1000;
        16'b0x1110x11110x10x : cnt0=17'h1000;
        16'b111110x11110x10x : cnt0=17'h2000;
        16'b0x0x0x111110x10x : cnt0=17'h800;
        16'b110x0x111110x10x : cnt0=17'h1000;
        16'b10x10x111110x10x : cnt0=17'h1000;
        16'b0x110x111110x10x : cnt0=17'h1000;
        16'b11110x111110x10x : cnt0=17'h2000;
        16'b10x0x1111110x10x : cnt0=17'h1000;
        16'b0x10x1111110x10x : cnt0=17'h1000;
        16'b1110x1111110x10x : cnt0=17'h2000;
        16'b0x0x11111110x10x : cnt0=17'h1000;
        16'b110x11111110x10x : cnt0=17'h2000;
        16'b10x111111110x10x : cnt0=17'h2000;
        16'b0x1111111110x10x : cnt0=17'h2000;
        16'b111111111110x10x : cnt0=17'h4000;
        16'b0x0x0x0x0x0x110x : cnt0=17'h200;
        16'b110x0x0x0x0x110x : cnt0=17'h400;
        16'b10x10x0x0x0x110x : cnt0=17'h400;
        16'b0x110x0x0x0x110x : cnt0=17'h400;
        16'b11110x0x0x0x110x : cnt0=17'h800;
        16'b10x0x10x0x0x110x : cnt0=17'h400;
        16'b0x10x10x0x0x110x : cnt0=17'h400;
        16'b1110x10x0x0x110x : cnt0=17'h800;
        16'b0x0x110x0x0x110x : cnt0=17'h400;
        16'b110x110x0x0x110x : cnt0=17'h800;
        16'b10x1110x0x0x110x : cnt0=17'h800;
        16'b0x11110x0x0x110x : cnt0=17'h800;
        16'b1111110x0x0x110x : cnt0=17'h1000;
        16'b10x0x0x10x0x110x : cnt0=17'h400;
        16'b0x10x0x10x0x110x : cnt0=17'h400;
        16'b1110x0x10x0x110x : cnt0=17'h800;
        16'b0x0x10x10x0x110x : cnt0=17'h400;
        16'b110x10x10x0x110x : cnt0=17'h800;
        16'b10x110x10x0x110x : cnt0=17'h800;
        16'b0x1110x10x0x110x : cnt0=17'h800;
        16'b111110x10x0x110x : cnt0=17'h1000;
        16'b0x0x0x110x0x110x : cnt0=17'h400;
        16'b110x0x110x0x110x : cnt0=17'h800;
        16'b10x10x110x0x110x : cnt0=17'h800;
        16'b0x110x110x0x110x : cnt0=17'h800;
        16'b11110x110x0x110x : cnt0=17'h1000;
        16'b10x0x1110x0x110x : cnt0=17'h800;
        16'b0x10x1110x0x110x : cnt0=17'h800;
        16'b1110x1110x0x110x : cnt0=17'h1000;
        16'b0x0x11110x0x110x : cnt0=17'h800;
        16'b110x11110x0x110x : cnt0=17'h1000;
        16'b10x111110x0x110x : cnt0=17'h1000;
        16'b0x1111110x0x110x : cnt0=17'h1000;
        16'b111111110x0x110x : cnt0=17'h2000;
        16'b10x0x0x0x10x110x : cnt0=17'h400;
        16'b0x10x0x0x10x110x : cnt0=17'h400;
        16'b1110x0x0x10x110x : cnt0=17'h800;
        16'b0x0x10x0x10x110x : cnt0=17'h400;
        16'b110x10x0x10x110x : cnt0=17'h800;
        16'b10x110x0x10x110x : cnt0=17'h800;
        16'b0x1110x0x10x110x : cnt0=17'h800;
        16'b111110x0x10x110x : cnt0=17'h1000;
        16'b0x0x0x10x10x110x : cnt0=17'h400;
        16'b110x0x10x10x110x : cnt0=17'h800;
        16'b10x10x10x10x110x : cnt0=17'h800;
        16'b0x110x10x10x110x : cnt0=17'h800;
        16'b11110x10x10x110x : cnt0=17'h1000;
        16'b10x0x110x10x110x : cnt0=17'h800;
        16'b0x10x110x10x110x : cnt0=17'h800;
        16'b1110x110x10x110x : cnt0=17'h1000;
        16'b0x0x1110x10x110x : cnt0=17'h800;
        16'b110x1110x10x110x : cnt0=17'h1000;
        16'b10x11110x10x110x : cnt0=17'h1000;
        16'b0x111110x10x110x : cnt0=17'h1000;
        16'b11111110x10x110x : cnt0=17'h2000;
        16'b0x0x0x0x110x110x : cnt0=17'h400;
        16'b110x0x0x110x110x : cnt0=17'h800;
        16'b10x10x0x110x110x : cnt0=17'h800;
        16'b0x110x0x110x110x : cnt0=17'h800;
        16'b11110x0x110x110x : cnt0=17'h1000;
        16'b10x0x10x110x110x : cnt0=17'h800;
        16'b0x10x10x110x110x : cnt0=17'h800;
        16'b1110x10x110x110x : cnt0=17'h1000;
        16'b0x0x110x110x110x : cnt0=17'h800;
        16'b110x110x110x110x : cnt0=17'h1000;
        16'b10x1110x110x110x : cnt0=17'h1000;
        16'b0x11110x110x110x : cnt0=17'h1000;
        16'b1111110x110x110x : cnt0=17'h2000;
        16'b10x0x0x1110x110x : cnt0=17'h800;
        16'b0x10x0x1110x110x : cnt0=17'h800;
        16'b1110x0x1110x110x : cnt0=17'h1000;
        16'b0x0x10x1110x110x : cnt0=17'h800;
        16'b110x10x1110x110x : cnt0=17'h1000;
        16'b10x110x1110x110x : cnt0=17'h1000;
        16'b0x1110x1110x110x : cnt0=17'h1000;
        16'b111110x1110x110x : cnt0=17'h2000;
        16'b0x0x0x11110x110x : cnt0=17'h800;
        16'b110x0x11110x110x : cnt0=17'h1000;
        16'b10x10x11110x110x : cnt0=17'h1000;
        16'b0x110x11110x110x : cnt0=17'h1000;
        16'b11110x11110x110x : cnt0=17'h2000;
        16'b10x0x111110x110x : cnt0=17'h1000;
        16'b0x10x111110x110x : cnt0=17'h1000;
        16'b1110x111110x110x : cnt0=17'h2000;
        16'b0x0x1111110x110x : cnt0=17'h1000;
        16'b110x1111110x110x : cnt0=17'h2000;
        16'b10x11111110x110x : cnt0=17'h2000;
        16'b0x111111110x110x : cnt0=17'h2000;
        16'b11111111110x110x : cnt0=17'h4000;
        16'b10x0x0x0x0x1110x : cnt0=17'h400;
        16'b0x10x0x0x0x1110x : cnt0=17'h400;
        16'b1110x0x0x0x1110x : cnt0=17'h800;
        16'b0x0x10x0x0x1110x : cnt0=17'h400;
        16'b110x10x0x0x1110x : cnt0=17'h800;
        16'b10x110x0x0x1110x : cnt0=17'h800;
        16'b0x1110x0x0x1110x : cnt0=17'h800;
        16'b111110x0x0x1110x : cnt0=17'h1000;
        16'b0x0x0x10x0x1110x : cnt0=17'h400;
        16'b110x0x10x0x1110x : cnt0=17'h800;
        16'b10x10x10x0x1110x : cnt0=17'h800;
        16'b0x110x10x0x1110x : cnt0=17'h800;
        16'b11110x10x0x1110x : cnt0=17'h1000;
        16'b10x0x110x0x1110x : cnt0=17'h800;
        16'b0x10x110x0x1110x : cnt0=17'h800;
        16'b1110x110x0x1110x : cnt0=17'h1000;
        16'b0x0x1110x0x1110x : cnt0=17'h800;
        16'b110x1110x0x1110x : cnt0=17'h1000;
        16'b10x11110x0x1110x : cnt0=17'h1000;
        16'b0x111110x0x1110x : cnt0=17'h1000;
        16'b11111110x0x1110x : cnt0=17'h2000;
        16'b0x0x0x0x10x1110x : cnt0=17'h400;
        16'b110x0x0x10x1110x : cnt0=17'h800;
        16'b10x10x0x10x1110x : cnt0=17'h800;
        16'b0x110x0x10x1110x : cnt0=17'h800;
        16'b11110x0x10x1110x : cnt0=17'h1000;
        16'b10x0x10x10x1110x : cnt0=17'h800;
        16'b0x10x10x10x1110x : cnt0=17'h800;
        16'b1110x10x10x1110x : cnt0=17'h1000;
        16'b0x0x110x10x1110x : cnt0=17'h800;
        16'b110x110x10x1110x : cnt0=17'h1000;
        16'b10x1110x10x1110x : cnt0=17'h1000;
        16'b0x11110x10x1110x : cnt0=17'h1000;
        16'b1111110x10x1110x : cnt0=17'h2000;
        16'b10x0x0x110x1110x : cnt0=17'h800;
        16'b0x10x0x110x1110x : cnt0=17'h800;
        16'b1110x0x110x1110x : cnt0=17'h1000;
        16'b0x0x10x110x1110x : cnt0=17'h800;
        16'b110x10x110x1110x : cnt0=17'h1000;
        16'b10x110x110x1110x : cnt0=17'h1000;
        16'b0x1110x110x1110x : cnt0=17'h1000;
        16'b111110x110x1110x : cnt0=17'h2000;
        16'b0x0x0x1110x1110x : cnt0=17'h800;
        16'b110x0x1110x1110x : cnt0=17'h1000;
        16'b10x10x1110x1110x : cnt0=17'h1000;
        16'b0x110x1110x1110x : cnt0=17'h1000;
        16'b11110x1110x1110x : cnt0=17'h2000;
        16'b10x0x11110x1110x : cnt0=17'h1000;
        16'b0x10x11110x1110x : cnt0=17'h1000;
        16'b1110x11110x1110x : cnt0=17'h2000;
        16'b0x0x111110x1110x : cnt0=17'h1000;
        16'b110x111110x1110x : cnt0=17'h2000;
        16'b10x1111110x1110x : cnt0=17'h2000;
        16'b0x11111110x1110x : cnt0=17'h2000;
        16'b1111111110x1110x : cnt0=17'h4000;
        16'b0x0x0x0x0x11110x : cnt0=17'h400;
        16'b110x0x0x0x11110x : cnt0=17'h800;
        16'b10x10x0x0x11110x : cnt0=17'h800;
        16'b0x110x0x0x11110x : cnt0=17'h800;
        16'b11110x0x0x11110x : cnt0=17'h1000;
        16'b10x0x10x0x11110x : cnt0=17'h800;
        16'b0x10x10x0x11110x : cnt0=17'h800;
        16'b1110x10x0x11110x : cnt0=17'h1000;
        16'b0x0x110x0x11110x : cnt0=17'h800;
        16'b110x110x0x11110x : cnt0=17'h1000;
        16'b10x1110x0x11110x : cnt0=17'h1000;
        16'b0x11110x0x11110x : cnt0=17'h1000;
        16'b1111110x0x11110x : cnt0=17'h2000;
        16'b10x0x0x10x11110x : cnt0=17'h800;
        16'b0x10x0x10x11110x : cnt0=17'h800;
        16'b1110x0x10x11110x : cnt0=17'h1000;
        16'b0x0x10x10x11110x : cnt0=17'h800;
        16'b110x10x10x11110x : cnt0=17'h1000;
        16'b10x110x10x11110x : cnt0=17'h1000;
        16'b0x1110x10x11110x : cnt0=17'h1000;
        16'b111110x10x11110x : cnt0=17'h2000;
        16'b0x0x0x110x11110x : cnt0=17'h800;
        16'b110x0x110x11110x : cnt0=17'h1000;
        16'b10x10x110x11110x : cnt0=17'h1000;
        16'b0x110x110x11110x : cnt0=17'h1000;
        16'b11110x110x11110x : cnt0=17'h2000;
        16'b10x0x1110x11110x : cnt0=17'h1000;
        16'b0x10x1110x11110x : cnt0=17'h1000;
        16'b1110x1110x11110x : cnt0=17'h2000;
        16'b0x0x11110x11110x : cnt0=17'h1000;
        16'b110x11110x11110x : cnt0=17'h2000;
        16'b10x111110x11110x : cnt0=17'h2000;
        16'b0x1111110x11110x : cnt0=17'h2000;
        16'b111111110x11110x : cnt0=17'h4000;
        16'b10x0x0x0x111110x : cnt0=17'h800;
        16'b0x10x0x0x111110x : cnt0=17'h800;
        16'b1110x0x0x111110x : cnt0=17'h1000;
        16'b0x0x10x0x111110x : cnt0=17'h800;
        16'b110x10x0x111110x : cnt0=17'h1000;
        16'b10x110x0x111110x : cnt0=17'h1000;
        16'b0x1110x0x111110x : cnt0=17'h1000;
        16'b111110x0x111110x : cnt0=17'h2000;
        16'b0x0x0x10x111110x : cnt0=17'h800;
        16'b110x0x10x111110x : cnt0=17'h1000;
        16'b10x10x10x111110x : cnt0=17'h1000;
        16'b0x110x10x111110x : cnt0=17'h1000;
        16'b11110x10x111110x : cnt0=17'h2000;
        16'b10x0x110x111110x : cnt0=17'h1000;
        16'b0x10x110x111110x : cnt0=17'h1000;
        16'b1110x110x111110x : cnt0=17'h2000;
        16'b0x0x1110x111110x : cnt0=17'h1000;
        16'b110x1110x111110x : cnt0=17'h2000;
        16'b10x11110x111110x : cnt0=17'h2000;
        16'b0x111110x111110x : cnt0=17'h2000;
        16'b11111110x111110x : cnt0=17'h4000;
        16'b0x0x0x0x1111110x : cnt0=17'h800;
        16'b110x0x0x1111110x : cnt0=17'h1000;
        16'b10x10x0x1111110x : cnt0=17'h1000;
        16'b0x110x0x1111110x : cnt0=17'h1000;
        16'b11110x0x1111110x : cnt0=17'h2000;
        16'b10x0x10x1111110x : cnt0=17'h1000;
        16'b0x10x10x1111110x : cnt0=17'h1000;
        16'b1110x10x1111110x : cnt0=17'h2000;
        16'b0x0x110x1111110x : cnt0=17'h1000;
        16'b110x110x1111110x : cnt0=17'h2000;
        16'b10x1110x1111110x : cnt0=17'h2000;
        16'b0x11110x1111110x : cnt0=17'h2000;
        16'b1111110x1111110x : cnt0=17'h4000;
        16'b10x0x0x11111110x : cnt0=17'h1000;
        16'b0x10x0x11111110x : cnt0=17'h1000;
        16'b1110x0x11111110x : cnt0=17'h2000;
        16'b0x0x10x11111110x : cnt0=17'h1000;
        16'b110x10x11111110x : cnt0=17'h2000;
        16'b10x110x11111110x : cnt0=17'h2000;
        16'b0x1110x11111110x : cnt0=17'h2000;
        16'b111110x11111110x : cnt0=17'h4000;
        16'b0x0x0x111111110x : cnt0=17'h1000;
        16'b110x0x111111110x : cnt0=17'h2000;
        16'b10x10x111111110x : cnt0=17'h2000;
        16'b0x110x111111110x : cnt0=17'h2000;
        16'b11110x111111110x : cnt0=17'h4000;
        16'b10x0x1111111110x : cnt0=17'h2000;
        16'b0x10x1111111110x : cnt0=17'h2000;
        16'b1110x1111111110x : cnt0=17'h4000;
        16'b0x0x11111111110x : cnt0=17'h2000;
        16'b110x11111111110x : cnt0=17'h4000;
        16'b10x111111111110x : cnt0=17'h4000;
        16'b0x1111111111110x : cnt0=17'h4000;
        16'b111111111111110x : cnt0=17'h8000;
        16'b0x0x0x0x0x0x0x10 : cnt0=17'h100;
        16'b110x0x0x0x0x0x10 : cnt0=17'h200;
        16'b10x10x0x0x0x0x10 : cnt0=17'h200;
        16'b0x110x0x0x0x0x10 : cnt0=17'h200;
        16'b11110x0x0x0x0x10 : cnt0=17'h400;
        16'b10x0x10x0x0x0x10 : cnt0=17'h200;
        16'b0x10x10x0x0x0x10 : cnt0=17'h200;
        16'b1110x10x0x0x0x10 : cnt0=17'h400;
        16'b0x0x110x0x0x0x10 : cnt0=17'h200;
        16'b110x110x0x0x0x10 : cnt0=17'h400;
        16'b10x1110x0x0x0x10 : cnt0=17'h400;
        16'b0x11110x0x0x0x10 : cnt0=17'h400;
        16'b1111110x0x0x0x10 : cnt0=17'h800;
        16'b10x0x0x10x0x0x10 : cnt0=17'h200;
        16'b0x10x0x10x0x0x10 : cnt0=17'h200;
        16'b1110x0x10x0x0x10 : cnt0=17'h400;
        16'b0x0x10x10x0x0x10 : cnt0=17'h200;
        16'b110x10x10x0x0x10 : cnt0=17'h400;
        16'b10x110x10x0x0x10 : cnt0=17'h400;
        16'b0x1110x10x0x0x10 : cnt0=17'h400;
        16'b111110x10x0x0x10 : cnt0=17'h800;
        16'b0x0x0x110x0x0x10 : cnt0=17'h200;
        16'b110x0x110x0x0x10 : cnt0=17'h400;
        16'b10x10x110x0x0x10 : cnt0=17'h400;
        16'b0x110x110x0x0x10 : cnt0=17'h400;
        16'b11110x110x0x0x10 : cnt0=17'h800;
        16'b10x0x1110x0x0x10 : cnt0=17'h400;
        16'b0x10x1110x0x0x10 : cnt0=17'h400;
        16'b1110x1110x0x0x10 : cnt0=17'h800;
        16'b0x0x11110x0x0x10 : cnt0=17'h400;
        16'b110x11110x0x0x10 : cnt0=17'h800;
        16'b10x111110x0x0x10 : cnt0=17'h800;
        16'b0x1111110x0x0x10 : cnt0=17'h800;
        16'b111111110x0x0x10 : cnt0=17'h1000;
        16'b10x0x0x0x10x0x10 : cnt0=17'h200;
        16'b0x10x0x0x10x0x10 : cnt0=17'h200;
        16'b1110x0x0x10x0x10 : cnt0=17'h400;
        16'b0x0x10x0x10x0x10 : cnt0=17'h200;
        16'b110x10x0x10x0x10 : cnt0=17'h400;
        16'b10x110x0x10x0x10 : cnt0=17'h400;
        16'b0x1110x0x10x0x10 : cnt0=17'h400;
        16'b111110x0x10x0x10 : cnt0=17'h800;
        16'b0x0x0x10x10x0x10 : cnt0=17'h200;
        16'b110x0x10x10x0x10 : cnt0=17'h400;
        16'b10x10x10x10x0x10 : cnt0=17'h400;
        16'b0x110x10x10x0x10 : cnt0=17'h400;
        16'b11110x10x10x0x10 : cnt0=17'h800;
        16'b10x0x110x10x0x10 : cnt0=17'h400;
        16'b0x10x110x10x0x10 : cnt0=17'h400;
        16'b1110x110x10x0x10 : cnt0=17'h800;
        16'b0x0x1110x10x0x10 : cnt0=17'h400;
        16'b110x1110x10x0x10 : cnt0=17'h800;
        16'b10x11110x10x0x10 : cnt0=17'h800;
        16'b0x111110x10x0x10 : cnt0=17'h800;
        16'b11111110x10x0x10 : cnt0=17'h1000;
        16'b0x0x0x0x110x0x10 : cnt0=17'h200;
        16'b110x0x0x110x0x10 : cnt0=17'h400;
        16'b10x10x0x110x0x10 : cnt0=17'h400;
        16'b0x110x0x110x0x10 : cnt0=17'h400;
        16'b11110x0x110x0x10 : cnt0=17'h800;
        16'b10x0x10x110x0x10 : cnt0=17'h400;
        16'b0x10x10x110x0x10 : cnt0=17'h400;
        16'b1110x10x110x0x10 : cnt0=17'h800;
        16'b0x0x110x110x0x10 : cnt0=17'h400;
        16'b110x110x110x0x10 : cnt0=17'h800;
        16'b10x1110x110x0x10 : cnt0=17'h800;
        16'b0x11110x110x0x10 : cnt0=17'h800;
        16'b1111110x110x0x10 : cnt0=17'h1000;
        16'b10x0x0x1110x0x10 : cnt0=17'h400;
        16'b0x10x0x1110x0x10 : cnt0=17'h400;
        16'b1110x0x1110x0x10 : cnt0=17'h800;
        16'b0x0x10x1110x0x10 : cnt0=17'h400;
        16'b110x10x1110x0x10 : cnt0=17'h800;
        16'b10x110x1110x0x10 : cnt0=17'h800;
        16'b0x1110x1110x0x10 : cnt0=17'h800;
        16'b111110x1110x0x10 : cnt0=17'h1000;
        16'b0x0x0x11110x0x10 : cnt0=17'h400;
        16'b110x0x11110x0x10 : cnt0=17'h800;
        16'b10x10x11110x0x10 : cnt0=17'h800;
        16'b0x110x11110x0x10 : cnt0=17'h800;
        16'b11110x11110x0x10 : cnt0=17'h1000;
        16'b10x0x111110x0x10 : cnt0=17'h800;
        16'b0x10x111110x0x10 : cnt0=17'h800;
        16'b1110x111110x0x10 : cnt0=17'h1000;
        16'b0x0x1111110x0x10 : cnt0=17'h800;
        16'b110x1111110x0x10 : cnt0=17'h1000;
        16'b10x11111110x0x10 : cnt0=17'h1000;
        16'b0x111111110x0x10 : cnt0=17'h1000;
        16'b11111111110x0x10 : cnt0=17'h2000;
        16'b10x0x0x0x0x10x10 : cnt0=17'h200;
        16'b0x10x0x0x0x10x10 : cnt0=17'h200;
        16'b1110x0x0x0x10x10 : cnt0=17'h400;
        16'b0x0x10x0x0x10x10 : cnt0=17'h200;
        16'b110x10x0x0x10x10 : cnt0=17'h400;
        16'b10x110x0x0x10x10 : cnt0=17'h400;
        16'b0x1110x0x0x10x10 : cnt0=17'h400;
        16'b111110x0x0x10x10 : cnt0=17'h800;
        16'b0x0x0x10x0x10x10 : cnt0=17'h200;
        16'b110x0x10x0x10x10 : cnt0=17'h400;
        16'b10x10x10x0x10x10 : cnt0=17'h400;
        16'b0x110x10x0x10x10 : cnt0=17'h400;
        16'b11110x10x0x10x10 : cnt0=17'h800;
        16'b10x0x110x0x10x10 : cnt0=17'h400;
        16'b0x10x110x0x10x10 : cnt0=17'h400;
        16'b1110x110x0x10x10 : cnt0=17'h800;
        16'b0x0x1110x0x10x10 : cnt0=17'h400;
        16'b110x1110x0x10x10 : cnt0=17'h800;
        16'b10x11110x0x10x10 : cnt0=17'h800;
        16'b0x111110x0x10x10 : cnt0=17'h800;
        16'b11111110x0x10x10 : cnt0=17'h1000;
        16'b0x0x0x0x10x10x10 : cnt0=17'h200;
        16'b110x0x0x10x10x10 : cnt0=17'h400;
        16'b10x10x0x10x10x10 : cnt0=17'h400;
        16'b0x110x0x10x10x10 : cnt0=17'h400;
        16'b11110x0x10x10x10 : cnt0=17'h800;
        16'b10x0x10x10x10x10 : cnt0=17'h400;
        16'b0x10x10x10x10x10 : cnt0=17'h400;
        16'b1110x10x10x10x10 : cnt0=17'h800;
        16'b0x0x110x10x10x10 : cnt0=17'h400;
        16'b110x110x10x10x10 : cnt0=17'h800;
        16'b10x1110x10x10x10 : cnt0=17'h800;
        16'b0x11110x10x10x10 : cnt0=17'h800;
        16'b1111110x10x10x10 : cnt0=17'h1000;
        16'b10x0x0x110x10x10 : cnt0=17'h400;
        16'b0x10x0x110x10x10 : cnt0=17'h400;
        16'b1110x0x110x10x10 : cnt0=17'h800;
        16'b0x0x10x110x10x10 : cnt0=17'h400;
        16'b110x10x110x10x10 : cnt0=17'h800;
        16'b10x110x110x10x10 : cnt0=17'h800;
        16'b0x1110x110x10x10 : cnt0=17'h800;
        16'b111110x110x10x10 : cnt0=17'h1000;
        16'b0x0x0x1110x10x10 : cnt0=17'h400;
        16'b110x0x1110x10x10 : cnt0=17'h800;
        16'b10x10x1110x10x10 : cnt0=17'h800;
        16'b0x110x1110x10x10 : cnt0=17'h800;
        16'b11110x1110x10x10 : cnt0=17'h1000;
        16'b10x0x11110x10x10 : cnt0=17'h800;
        16'b0x10x11110x10x10 : cnt0=17'h800;
        16'b1110x11110x10x10 : cnt0=17'h1000;
        16'b0x0x111110x10x10 : cnt0=17'h800;
        16'b110x111110x10x10 : cnt0=17'h1000;
        16'b10x1111110x10x10 : cnt0=17'h1000;
        16'b0x11111110x10x10 : cnt0=17'h1000;
        16'b1111111110x10x10 : cnt0=17'h2000;
        16'b0x0x0x0x0x110x10 : cnt0=17'h200;
        16'b110x0x0x0x110x10 : cnt0=17'h400;
        16'b10x10x0x0x110x10 : cnt0=17'h400;
        16'b0x110x0x0x110x10 : cnt0=17'h400;
        16'b11110x0x0x110x10 : cnt0=17'h800;
        16'b10x0x10x0x110x10 : cnt0=17'h400;
        16'b0x10x10x0x110x10 : cnt0=17'h400;
        16'b1110x10x0x110x10 : cnt0=17'h800;
        16'b0x0x110x0x110x10 : cnt0=17'h400;
        16'b110x110x0x110x10 : cnt0=17'h800;
        16'b10x1110x0x110x10 : cnt0=17'h800;
        16'b0x11110x0x110x10 : cnt0=17'h800;
        16'b1111110x0x110x10 : cnt0=17'h1000;
        16'b10x0x0x10x110x10 : cnt0=17'h400;
        16'b0x10x0x10x110x10 : cnt0=17'h400;
        16'b1110x0x10x110x10 : cnt0=17'h800;
        16'b0x0x10x10x110x10 : cnt0=17'h400;
        16'b110x10x10x110x10 : cnt0=17'h800;
        16'b10x110x10x110x10 : cnt0=17'h800;
        16'b0x1110x10x110x10 : cnt0=17'h800;
        16'b111110x10x110x10 : cnt0=17'h1000;
        16'b0x0x0x110x110x10 : cnt0=17'h400;
        16'b110x0x110x110x10 : cnt0=17'h800;
        16'b10x10x110x110x10 : cnt0=17'h800;
        16'b0x110x110x110x10 : cnt0=17'h800;
        16'b11110x110x110x10 : cnt0=17'h1000;
        16'b10x0x1110x110x10 : cnt0=17'h800;
        16'b0x10x1110x110x10 : cnt0=17'h800;
        16'b1110x1110x110x10 : cnt0=17'h1000;
        16'b0x0x11110x110x10 : cnt0=17'h800;
        16'b110x11110x110x10 : cnt0=17'h1000;
        16'b10x111110x110x10 : cnt0=17'h1000;
        16'b0x1111110x110x10 : cnt0=17'h1000;
        16'b111111110x110x10 : cnt0=17'h2000;
        16'b10x0x0x0x1110x10 : cnt0=17'h400;
        16'b0x10x0x0x1110x10 : cnt0=17'h400;
        16'b1110x0x0x1110x10 : cnt0=17'h800;
        16'b0x0x10x0x1110x10 : cnt0=17'h400;
        16'b110x10x0x1110x10 : cnt0=17'h800;
        16'b10x110x0x1110x10 : cnt0=17'h800;
        16'b0x1110x0x1110x10 : cnt0=17'h800;
        16'b111110x0x1110x10 : cnt0=17'h1000;
        16'b0x0x0x10x1110x10 : cnt0=17'h400;
        16'b110x0x10x1110x10 : cnt0=17'h800;
        16'b10x10x10x1110x10 : cnt0=17'h800;
        16'b0x110x10x1110x10 : cnt0=17'h800;
        16'b11110x10x1110x10 : cnt0=17'h1000;
        16'b10x0x110x1110x10 : cnt0=17'h800;
        16'b0x10x110x1110x10 : cnt0=17'h800;
        16'b1110x110x1110x10 : cnt0=17'h1000;
        16'b0x0x1110x1110x10 : cnt0=17'h800;
        16'b110x1110x1110x10 : cnt0=17'h1000;
        16'b10x11110x1110x10 : cnt0=17'h1000;
        16'b0x111110x1110x10 : cnt0=17'h1000;
        16'b11111110x1110x10 : cnt0=17'h2000;
        16'b0x0x0x0x11110x10 : cnt0=17'h400;
        16'b110x0x0x11110x10 : cnt0=17'h800;
        16'b10x10x0x11110x10 : cnt0=17'h800;
        16'b0x110x0x11110x10 : cnt0=17'h800;
        16'b11110x0x11110x10 : cnt0=17'h1000;
        16'b10x0x10x11110x10 : cnt0=17'h800;
        16'b0x10x10x11110x10 : cnt0=17'h800;
        16'b1110x10x11110x10 : cnt0=17'h1000;
        16'b0x0x110x11110x10 : cnt0=17'h800;
        16'b110x110x11110x10 : cnt0=17'h1000;
        16'b10x1110x11110x10 : cnt0=17'h1000;
        16'b0x11110x11110x10 : cnt0=17'h1000;
        16'b1111110x11110x10 : cnt0=17'h2000;
        16'b10x0x0x111110x10 : cnt0=17'h800;
        16'b0x10x0x111110x10 : cnt0=17'h800;
        16'b1110x0x111110x10 : cnt0=17'h1000;
        16'b0x0x10x111110x10 : cnt0=17'h800;
        16'b110x10x111110x10 : cnt0=17'h1000;
        16'b10x110x111110x10 : cnt0=17'h1000;
        16'b0x1110x111110x10 : cnt0=17'h1000;
        16'b111110x111110x10 : cnt0=17'h2000;
        16'b0x0x0x1111110x10 : cnt0=17'h800;
        16'b110x0x1111110x10 : cnt0=17'h1000;
        16'b10x10x1111110x10 : cnt0=17'h1000;
        16'b0x110x1111110x10 : cnt0=17'h1000;
        16'b11110x1111110x10 : cnt0=17'h2000;
        16'b10x0x11111110x10 : cnt0=17'h1000;
        16'b0x10x11111110x10 : cnt0=17'h1000;
        16'b1110x11111110x10 : cnt0=17'h2000;
        16'b0x0x111111110x10 : cnt0=17'h1000;
        16'b110x111111110x10 : cnt0=17'h2000;
        16'b10x1111111110x10 : cnt0=17'h2000;
        16'b0x11111111110x10 : cnt0=17'h2000;
        16'b1111111111110x10 : cnt0=17'h4000;
        16'b10x0x0x0x0x0x110 : cnt0=17'h200;
        16'b0x10x0x0x0x0x110 : cnt0=17'h200;
        16'b1110x0x0x0x0x110 : cnt0=17'h400;
        16'b0x0x10x0x0x0x110 : cnt0=17'h200;
        16'b110x10x0x0x0x110 : cnt0=17'h400;
        16'b10x110x0x0x0x110 : cnt0=17'h400;
        16'b0x1110x0x0x0x110 : cnt0=17'h400;
        16'b111110x0x0x0x110 : cnt0=17'h800;
        16'b0x0x0x10x0x0x110 : cnt0=17'h200;
        16'b110x0x10x0x0x110 : cnt0=17'h400;
        16'b10x10x10x0x0x110 : cnt0=17'h400;
        16'b0x110x10x0x0x110 : cnt0=17'h400;
        16'b11110x10x0x0x110 : cnt0=17'h800;
        16'b10x0x110x0x0x110 : cnt0=17'h400;
        16'b0x10x110x0x0x110 : cnt0=17'h400;
        16'b1110x110x0x0x110 : cnt0=17'h800;
        16'b0x0x1110x0x0x110 : cnt0=17'h400;
        16'b110x1110x0x0x110 : cnt0=17'h800;
        16'b10x11110x0x0x110 : cnt0=17'h800;
        16'b0x111110x0x0x110 : cnt0=17'h800;
        16'b11111110x0x0x110 : cnt0=17'h1000;
        16'b0x0x0x0x10x0x110 : cnt0=17'h200;
        16'b110x0x0x10x0x110 : cnt0=17'h400;
        16'b10x10x0x10x0x110 : cnt0=17'h400;
        16'b0x110x0x10x0x110 : cnt0=17'h400;
        16'b11110x0x10x0x110 : cnt0=17'h800;
        16'b10x0x10x10x0x110 : cnt0=17'h400;
        16'b0x10x10x10x0x110 : cnt0=17'h400;
        16'b1110x10x10x0x110 : cnt0=17'h800;
        16'b0x0x110x10x0x110 : cnt0=17'h400;
        16'b110x110x10x0x110 : cnt0=17'h800;
        16'b10x1110x10x0x110 : cnt0=17'h800;
        16'b0x11110x10x0x110 : cnt0=17'h800;
        16'b1111110x10x0x110 : cnt0=17'h1000;
        16'b10x0x0x110x0x110 : cnt0=17'h400;
        16'b0x10x0x110x0x110 : cnt0=17'h400;
        16'b1110x0x110x0x110 : cnt0=17'h800;
        16'b0x0x10x110x0x110 : cnt0=17'h400;
        16'b110x10x110x0x110 : cnt0=17'h800;
        16'b10x110x110x0x110 : cnt0=17'h800;
        16'b0x1110x110x0x110 : cnt0=17'h800;
        16'b111110x110x0x110 : cnt0=17'h1000;
        16'b0x0x0x1110x0x110 : cnt0=17'h400;
        16'b110x0x1110x0x110 : cnt0=17'h800;
        16'b10x10x1110x0x110 : cnt0=17'h800;
        16'b0x110x1110x0x110 : cnt0=17'h800;
        16'b11110x1110x0x110 : cnt0=17'h1000;
        16'b10x0x11110x0x110 : cnt0=17'h800;
        16'b0x10x11110x0x110 : cnt0=17'h800;
        16'b1110x11110x0x110 : cnt0=17'h1000;
        16'b0x0x111110x0x110 : cnt0=17'h800;
        16'b110x111110x0x110 : cnt0=17'h1000;
        16'b10x1111110x0x110 : cnt0=17'h1000;
        16'b0x11111110x0x110 : cnt0=17'h1000;
        16'b1111111110x0x110 : cnt0=17'h2000;
        16'b0x0x0x0x0x10x110 : cnt0=17'h200;
        16'b110x0x0x0x10x110 : cnt0=17'h400;
        16'b10x10x0x0x10x110 : cnt0=17'h400;
        16'b0x110x0x0x10x110 : cnt0=17'h400;
        16'b11110x0x0x10x110 : cnt0=17'h800;
        16'b10x0x10x0x10x110 : cnt0=17'h400;
        16'b0x10x10x0x10x110 : cnt0=17'h400;
        16'b1110x10x0x10x110 : cnt0=17'h800;
        16'b0x0x110x0x10x110 : cnt0=17'h400;
        16'b110x110x0x10x110 : cnt0=17'h800;
        16'b10x1110x0x10x110 : cnt0=17'h800;
        16'b0x11110x0x10x110 : cnt0=17'h800;
        16'b1111110x0x10x110 : cnt0=17'h1000;
        16'b10x0x0x10x10x110 : cnt0=17'h400;
        16'b0x10x0x10x10x110 : cnt0=17'h400;
        16'b1110x0x10x10x110 : cnt0=17'h800;
        16'b0x0x10x10x10x110 : cnt0=17'h400;
        16'b110x10x10x10x110 : cnt0=17'h800;
        16'b10x110x10x10x110 : cnt0=17'h800;
        16'b0x1110x10x10x110 : cnt0=17'h800;
        16'b111110x10x10x110 : cnt0=17'h1000;
        16'b0x0x0x110x10x110 : cnt0=17'h400;
        16'b110x0x110x10x110 : cnt0=17'h800;
        16'b10x10x110x10x110 : cnt0=17'h800;
        16'b0x110x110x10x110 : cnt0=17'h800;
        16'b11110x110x10x110 : cnt0=17'h1000;
        16'b10x0x1110x10x110 : cnt0=17'h800;
        16'b0x10x1110x10x110 : cnt0=17'h800;
        16'b1110x1110x10x110 : cnt0=17'h1000;
        16'b0x0x11110x10x110 : cnt0=17'h800;
        16'b110x11110x10x110 : cnt0=17'h1000;
        16'b10x111110x10x110 : cnt0=17'h1000;
        16'b0x1111110x10x110 : cnt0=17'h1000;
        16'b111111110x10x110 : cnt0=17'h2000;
        16'b10x0x0x0x110x110 : cnt0=17'h400;
        16'b0x10x0x0x110x110 : cnt0=17'h400;
        16'b1110x0x0x110x110 : cnt0=17'h800;
        16'b0x0x10x0x110x110 : cnt0=17'h400;
        16'b110x10x0x110x110 : cnt0=17'h800;
        16'b10x110x0x110x110 : cnt0=17'h800;
        16'b0x1110x0x110x110 : cnt0=17'h800;
        16'b111110x0x110x110 : cnt0=17'h1000;
        16'b0x0x0x10x110x110 : cnt0=17'h400;
        16'b110x0x10x110x110 : cnt0=17'h800;
        16'b10x10x10x110x110 : cnt0=17'h800;
        16'b0x110x10x110x110 : cnt0=17'h800;
        16'b11110x10x110x110 : cnt0=17'h1000;
        16'b10x0x110x110x110 : cnt0=17'h800;
        16'b0x10x110x110x110 : cnt0=17'h800;
        16'b1110x110x110x110 : cnt0=17'h1000;
        16'b0x0x1110x110x110 : cnt0=17'h800;
        16'b110x1110x110x110 : cnt0=17'h1000;
        16'b10x11110x110x110 : cnt0=17'h1000;
        16'b0x111110x110x110 : cnt0=17'h1000;
        16'b11111110x110x110 : cnt0=17'h2000;
        16'b0x0x0x0x1110x110 : cnt0=17'h400;
        16'b110x0x0x1110x110 : cnt0=17'h800;
        16'b10x10x0x1110x110 : cnt0=17'h800;
        16'b0x110x0x1110x110 : cnt0=17'h800;
        16'b11110x0x1110x110 : cnt0=17'h1000;
        16'b10x0x10x1110x110 : cnt0=17'h800;
        16'b0x10x10x1110x110 : cnt0=17'h800;
        16'b1110x10x1110x110 : cnt0=17'h1000;
        16'b0x0x110x1110x110 : cnt0=17'h800;
        16'b110x110x1110x110 : cnt0=17'h1000;
        16'b10x1110x1110x110 : cnt0=17'h1000;
        16'b0x11110x1110x110 : cnt0=17'h1000;
        16'b1111110x1110x110 : cnt0=17'h2000;
        16'b10x0x0x11110x110 : cnt0=17'h800;
        16'b0x10x0x11110x110 : cnt0=17'h800;
        16'b1110x0x11110x110 : cnt0=17'h1000;
        16'b0x0x10x11110x110 : cnt0=17'h800;
        16'b110x10x11110x110 : cnt0=17'h1000;
        16'b10x110x11110x110 : cnt0=17'h1000;
        16'b0x1110x11110x110 : cnt0=17'h1000;
        16'b111110x11110x110 : cnt0=17'h2000;
        16'b0x0x0x111110x110 : cnt0=17'h800;
        16'b110x0x111110x110 : cnt0=17'h1000;
        16'b10x10x111110x110 : cnt0=17'h1000;
        16'b0x110x111110x110 : cnt0=17'h1000;
        16'b11110x111110x110 : cnt0=17'h2000;
        16'b10x0x1111110x110 : cnt0=17'h1000;
        16'b0x10x1111110x110 : cnt0=17'h1000;
        16'b1110x1111110x110 : cnt0=17'h2000;
        16'b0x0x11111110x110 : cnt0=17'h1000;
        16'b110x11111110x110 : cnt0=17'h2000;
        16'b10x111111110x110 : cnt0=17'h2000;
        16'b0x1111111110x110 : cnt0=17'h2000;
        16'b111111111110x110 : cnt0=17'h4000;
        16'b0x0x0x0x0x0x1110 : cnt0=17'h200;
        16'b110x0x0x0x0x1110 : cnt0=17'h400;
        16'b10x10x0x0x0x1110 : cnt0=17'h400;
        16'b0x110x0x0x0x1110 : cnt0=17'h400;
        16'b11110x0x0x0x1110 : cnt0=17'h800;
        16'b10x0x10x0x0x1110 : cnt0=17'h400;
        16'b0x10x10x0x0x1110 : cnt0=17'h400;
        16'b1110x10x0x0x1110 : cnt0=17'h800;
        16'b0x0x110x0x0x1110 : cnt0=17'h400;
        16'b110x110x0x0x1110 : cnt0=17'h800;
        16'b10x1110x0x0x1110 : cnt0=17'h800;
        16'b0x11110x0x0x1110 : cnt0=17'h800;
        16'b1111110x0x0x1110 : cnt0=17'h1000;
        16'b10x0x0x10x0x1110 : cnt0=17'h400;
        16'b0x10x0x10x0x1110 : cnt0=17'h400;
        16'b1110x0x10x0x1110 : cnt0=17'h800;
        16'b0x0x10x10x0x1110 : cnt0=17'h400;
        16'b110x10x10x0x1110 : cnt0=17'h800;
        16'b10x110x10x0x1110 : cnt0=17'h800;
        16'b0x1110x10x0x1110 : cnt0=17'h800;
        16'b111110x10x0x1110 : cnt0=17'h1000;
        16'b0x0x0x110x0x1110 : cnt0=17'h400;
        16'b110x0x110x0x1110 : cnt0=17'h800;
        16'b10x10x110x0x1110 : cnt0=17'h800;
        16'b0x110x110x0x1110 : cnt0=17'h800;
        16'b11110x110x0x1110 : cnt0=17'h1000;
        16'b10x0x1110x0x1110 : cnt0=17'h800;
        16'b0x10x1110x0x1110 : cnt0=17'h800;
        16'b1110x1110x0x1110 : cnt0=17'h1000;
        16'b0x0x11110x0x1110 : cnt0=17'h800;
        16'b110x11110x0x1110 : cnt0=17'h1000;
        16'b10x111110x0x1110 : cnt0=17'h1000;
        16'b0x1111110x0x1110 : cnt0=17'h1000;
        16'b111111110x0x1110 : cnt0=17'h2000;
        16'b10x0x0x0x10x1110 : cnt0=17'h400;
        16'b0x10x0x0x10x1110 : cnt0=17'h400;
        16'b1110x0x0x10x1110 : cnt0=17'h800;
        16'b0x0x10x0x10x1110 : cnt0=17'h400;
        16'b110x10x0x10x1110 : cnt0=17'h800;
        16'b10x110x0x10x1110 : cnt0=17'h800;
        16'b0x1110x0x10x1110 : cnt0=17'h800;
        16'b111110x0x10x1110 : cnt0=17'h1000;
        16'b0x0x0x10x10x1110 : cnt0=17'h400;
        16'b110x0x10x10x1110 : cnt0=17'h800;
        16'b10x10x10x10x1110 : cnt0=17'h800;
        16'b0x110x10x10x1110 : cnt0=17'h800;
        16'b11110x10x10x1110 : cnt0=17'h1000;
        16'b10x0x110x10x1110 : cnt0=17'h800;
        16'b0x10x110x10x1110 : cnt0=17'h800;
        16'b1110x110x10x1110 : cnt0=17'h1000;
        16'b0x0x1110x10x1110 : cnt0=17'h800;
        16'b110x1110x10x1110 : cnt0=17'h1000;
        16'b10x11110x10x1110 : cnt0=17'h1000;
        16'b0x111110x10x1110 : cnt0=17'h1000;
        16'b11111110x10x1110 : cnt0=17'h2000;
        16'b0x0x0x0x110x1110 : cnt0=17'h400;
        16'b110x0x0x110x1110 : cnt0=17'h800;
        16'b10x10x0x110x1110 : cnt0=17'h800;
        16'b0x110x0x110x1110 : cnt0=17'h800;
        16'b11110x0x110x1110 : cnt0=17'h1000;
        16'b10x0x10x110x1110 : cnt0=17'h800;
        16'b0x10x10x110x1110 : cnt0=17'h800;
        16'b1110x10x110x1110 : cnt0=17'h1000;
        16'b0x0x110x110x1110 : cnt0=17'h800;
        16'b110x110x110x1110 : cnt0=17'h1000;
        16'b10x1110x110x1110 : cnt0=17'h1000;
        16'b0x11110x110x1110 : cnt0=17'h1000;
        16'b1111110x110x1110 : cnt0=17'h2000;
        16'b10x0x0x1110x1110 : cnt0=17'h800;
        16'b0x10x0x1110x1110 : cnt0=17'h800;
        16'b1110x0x1110x1110 : cnt0=17'h1000;
        16'b0x0x10x1110x1110 : cnt0=17'h800;
        16'b110x10x1110x1110 : cnt0=17'h1000;
        16'b10x110x1110x1110 : cnt0=17'h1000;
        16'b0x1110x1110x1110 : cnt0=17'h1000;
        16'b111110x1110x1110 : cnt0=17'h2000;
        16'b0x0x0x11110x1110 : cnt0=17'h800;
        16'b110x0x11110x1110 : cnt0=17'h1000;
        16'b10x10x11110x1110 : cnt0=17'h1000;
        16'b0x110x11110x1110 : cnt0=17'h1000;
        16'b11110x11110x1110 : cnt0=17'h2000;
        16'b10x0x111110x1110 : cnt0=17'h1000;
        16'b0x10x111110x1110 : cnt0=17'h1000;
        16'b1110x111110x1110 : cnt0=17'h2000;
        16'b0x0x1111110x1110 : cnt0=17'h1000;
        16'b110x1111110x1110 : cnt0=17'h2000;
        16'b10x11111110x1110 : cnt0=17'h2000;
        16'b0x111111110x1110 : cnt0=17'h2000;
        16'b11111111110x1110 : cnt0=17'h4000;
        16'b10x0x0x0x0x11110 : cnt0=17'h400;
        16'b0x10x0x0x0x11110 : cnt0=17'h400;
        16'b1110x0x0x0x11110 : cnt0=17'h800;
        16'b0x0x10x0x0x11110 : cnt0=17'h400;
        16'b110x10x0x0x11110 : cnt0=17'h800;
        16'b10x110x0x0x11110 : cnt0=17'h800;
        16'b0x1110x0x0x11110 : cnt0=17'h800;
        16'b111110x0x0x11110 : cnt0=17'h1000;
        16'b0x0x0x10x0x11110 : cnt0=17'h400;
        16'b110x0x10x0x11110 : cnt0=17'h800;
        16'b10x10x10x0x11110 : cnt0=17'h800;
        16'b0x110x10x0x11110 : cnt0=17'h800;
        16'b11110x10x0x11110 : cnt0=17'h1000;
        16'b10x0x110x0x11110 : cnt0=17'h800;
        16'b0x10x110x0x11110 : cnt0=17'h800;
        16'b1110x110x0x11110 : cnt0=17'h1000;
        16'b0x0x1110x0x11110 : cnt0=17'h800;
        16'b110x1110x0x11110 : cnt0=17'h1000;
        16'b10x11110x0x11110 : cnt0=17'h1000;
        16'b0x111110x0x11110 : cnt0=17'h1000;
        16'b11111110x0x11110 : cnt0=17'h2000;
        16'b0x0x0x0x10x11110 : cnt0=17'h400;
        16'b110x0x0x10x11110 : cnt0=17'h800;
        16'b10x10x0x10x11110 : cnt0=17'h800;
        16'b0x110x0x10x11110 : cnt0=17'h800;
        16'b11110x0x10x11110 : cnt0=17'h1000;
        16'b10x0x10x10x11110 : cnt0=17'h800;
        16'b0x10x10x10x11110 : cnt0=17'h800;
        16'b1110x10x10x11110 : cnt0=17'h1000;
        16'b0x0x110x10x11110 : cnt0=17'h800;
        16'b110x110x10x11110 : cnt0=17'h1000;
        16'b10x1110x10x11110 : cnt0=17'h1000;
        16'b0x11110x10x11110 : cnt0=17'h1000;
        16'b1111110x10x11110 : cnt0=17'h2000;
        16'b10x0x0x110x11110 : cnt0=17'h800;
        16'b0x10x0x110x11110 : cnt0=17'h800;
        16'b1110x0x110x11110 : cnt0=17'h1000;
        16'b0x0x10x110x11110 : cnt0=17'h800;
        16'b110x10x110x11110 : cnt0=17'h1000;
        16'b10x110x110x11110 : cnt0=17'h1000;
        16'b0x1110x110x11110 : cnt0=17'h1000;
        16'b111110x110x11110 : cnt0=17'h2000;
        16'b0x0x0x1110x11110 : cnt0=17'h800;
        16'b110x0x1110x11110 : cnt0=17'h1000;
        16'b10x10x1110x11110 : cnt0=17'h1000;
        16'b0x110x1110x11110 : cnt0=17'h1000;
        16'b11110x1110x11110 : cnt0=17'h2000;
        16'b10x0x11110x11110 : cnt0=17'h1000;
        16'b0x10x11110x11110 : cnt0=17'h1000;
        16'b1110x11110x11110 : cnt0=17'h2000;
        16'b0x0x111110x11110 : cnt0=17'h1000;
        16'b110x111110x11110 : cnt0=17'h2000;
        16'b10x1111110x11110 : cnt0=17'h2000;
        16'b0x11111110x11110 : cnt0=17'h2000;
        16'b1111111110x11110 : cnt0=17'h4000;
        16'b0x0x0x0x0x111110 : cnt0=17'h400;
        16'b110x0x0x0x111110 : cnt0=17'h800;
        16'b10x10x0x0x111110 : cnt0=17'h800;
        16'b0x110x0x0x111110 : cnt0=17'h800;
        16'b11110x0x0x111110 : cnt0=17'h1000;
        16'b10x0x10x0x111110 : cnt0=17'h800;
        16'b0x10x10x0x111110 : cnt0=17'h800;
        16'b1110x10x0x111110 : cnt0=17'h1000;
        16'b0x0x110x0x111110 : cnt0=17'h800;
        16'b110x110x0x111110 : cnt0=17'h1000;
        16'b10x1110x0x111110 : cnt0=17'h1000;
        16'b0x11110x0x111110 : cnt0=17'h1000;
        16'b1111110x0x111110 : cnt0=17'h2000;
        16'b10x0x0x10x111110 : cnt0=17'h800;
        16'b0x10x0x10x111110 : cnt0=17'h800;
        16'b1110x0x10x111110 : cnt0=17'h1000;
        16'b0x0x10x10x111110 : cnt0=17'h800;
        16'b110x10x10x111110 : cnt0=17'h1000;
        16'b10x110x10x111110 : cnt0=17'h1000;
        16'b0x1110x10x111110 : cnt0=17'h1000;
        16'b111110x10x111110 : cnt0=17'h2000;
        16'b0x0x0x110x111110 : cnt0=17'h800;
        16'b110x0x110x111110 : cnt0=17'h1000;
        16'b10x10x110x111110 : cnt0=17'h1000;
        16'b0x110x110x111110 : cnt0=17'h1000;
        16'b11110x110x111110 : cnt0=17'h2000;
        16'b10x0x1110x111110 : cnt0=17'h1000;
        16'b0x10x1110x111110 : cnt0=17'h1000;
        16'b1110x1110x111110 : cnt0=17'h2000;
        16'b0x0x11110x111110 : cnt0=17'h1000;
        16'b110x11110x111110 : cnt0=17'h2000;
        16'b10x111110x111110 : cnt0=17'h2000;
        16'b0x1111110x111110 : cnt0=17'h2000;
        16'b111111110x111110 : cnt0=17'h4000;
        16'b10x0x0x0x1111110 : cnt0=17'h800;
        16'b0x10x0x0x1111110 : cnt0=17'h800;
        16'b1110x0x0x1111110 : cnt0=17'h1000;
        16'b0x0x10x0x1111110 : cnt0=17'h800;
        16'b110x10x0x1111110 : cnt0=17'h1000;
        16'b10x110x0x1111110 : cnt0=17'h1000;
        16'b0x1110x0x1111110 : cnt0=17'h1000;
        16'b111110x0x1111110 : cnt0=17'h2000;
        16'b0x0x0x10x1111110 : cnt0=17'h800;
        16'b110x0x10x1111110 : cnt0=17'h1000;
        16'b10x10x10x1111110 : cnt0=17'h1000;
        16'b0x110x10x1111110 : cnt0=17'h1000;
        16'b11110x10x1111110 : cnt0=17'h2000;
        16'b10x0x110x1111110 : cnt0=17'h1000;
        16'b0x10x110x1111110 : cnt0=17'h1000;
        16'b1110x110x1111110 : cnt0=17'h2000;
        16'b0x0x1110x1111110 : cnt0=17'h1000;
        16'b110x1110x1111110 : cnt0=17'h2000;
        16'b10x11110x1111110 : cnt0=17'h2000;
        16'b0x111110x1111110 : cnt0=17'h2000;
        16'b11111110x1111110 : cnt0=17'h4000;
        16'b0x0x0x0x11111110 : cnt0=17'h800;
        16'b110x0x0x11111110 : cnt0=17'h1000;
        16'b10x10x0x11111110 : cnt0=17'h1000;
        16'b0x110x0x11111110 : cnt0=17'h1000;
        16'b11110x0x11111110 : cnt0=17'h2000;
        16'b10x0x10x11111110 : cnt0=17'h1000;
        16'b0x10x10x11111110 : cnt0=17'h1000;
        16'b1110x10x11111110 : cnt0=17'h2000;
        16'b0x0x110x11111110 : cnt0=17'h1000;
        16'b110x110x11111110 : cnt0=17'h2000;
        16'b10x1110x11111110 : cnt0=17'h2000;
        16'b0x11110x11111110 : cnt0=17'h2000;
        16'b1111110x11111110 : cnt0=17'h4000;
        16'b10x0x0x111111110 : cnt0=17'h1000;
        16'b0x10x0x111111110 : cnt0=17'h1000;
        16'b1110x0x111111110 : cnt0=17'h2000;
        16'b0x0x10x111111110 : cnt0=17'h1000;
        16'b110x10x111111110 : cnt0=17'h2000;
        16'b10x110x111111110 : cnt0=17'h2000;
        16'b0x1110x111111110 : cnt0=17'h2000;
        16'b111110x111111110 : cnt0=17'h4000;
        16'b0x0x0x1111111110 : cnt0=17'h1000;
        16'b110x0x1111111110 : cnt0=17'h2000;
        16'b10x10x1111111110 : cnt0=17'h2000;
        16'b0x110x1111111110 : cnt0=17'h2000;
        16'b11110x1111111110 : cnt0=17'h4000;
        16'b10x0x11111111110 : cnt0=17'h2000;
        16'b0x10x11111111110 : cnt0=17'h2000;
        16'b1110x11111111110 : cnt0=17'h4000;
        16'b0x0x111111111110 : cnt0=17'h2000;
        16'b110x111111111110 : cnt0=17'h4000;
        16'b10x1111111111110 : cnt0=17'h4000;
        16'b0x11111111111110 : cnt0=17'h4000;
        16'b1111111111111110 : cnt0=17'h8000;
        16'b10x0x0x0x0x0x0x1 : cnt0=17'h200;
        16'b0x10x0x0x0x0x0x1 : cnt0=17'h200;
        16'b1110x0x0x0x0x0x1 : cnt0=17'h400;
        16'b0x0x10x0x0x0x0x1 : cnt0=17'h200;
        16'b110x10x0x0x0x0x1 : cnt0=17'h400;
        16'b10x110x0x0x0x0x1 : cnt0=17'h400;
        16'b0x1110x0x0x0x0x1 : cnt0=17'h400;
        16'b111110x0x0x0x0x1 : cnt0=17'h800;
        16'b0x0x0x10x0x0x0x1 : cnt0=17'h200;
        16'b110x0x10x0x0x0x1 : cnt0=17'h400;
        16'b10x10x10x0x0x0x1 : cnt0=17'h400;
        16'b0x110x10x0x0x0x1 : cnt0=17'h400;
        16'b11110x10x0x0x0x1 : cnt0=17'h800;
        16'b10x0x110x0x0x0x1 : cnt0=17'h400;
        16'b0x10x110x0x0x0x1 : cnt0=17'h400;
        16'b1110x110x0x0x0x1 : cnt0=17'h800;
        16'b0x0x1110x0x0x0x1 : cnt0=17'h400;
        16'b110x1110x0x0x0x1 : cnt0=17'h800;
        16'b10x11110x0x0x0x1 : cnt0=17'h800;
        16'b0x111110x0x0x0x1 : cnt0=17'h800;
        16'b11111110x0x0x0x1 : cnt0=17'h1000;
        16'b0x0x0x0x10x0x0x1 : cnt0=17'h200;
        16'b110x0x0x10x0x0x1 : cnt0=17'h400;
        16'b10x10x0x10x0x0x1 : cnt0=17'h400;
        16'b0x110x0x10x0x0x1 : cnt0=17'h400;
        16'b11110x0x10x0x0x1 : cnt0=17'h800;
        16'b10x0x10x10x0x0x1 : cnt0=17'h400;
        16'b0x10x10x10x0x0x1 : cnt0=17'h400;
        16'b1110x10x10x0x0x1 : cnt0=17'h800;
        16'b0x0x110x10x0x0x1 : cnt0=17'h400;
        16'b110x110x10x0x0x1 : cnt0=17'h800;
        16'b10x1110x10x0x0x1 : cnt0=17'h800;
        16'b0x11110x10x0x0x1 : cnt0=17'h800;
        16'b1111110x10x0x0x1 : cnt0=17'h1000;
        16'b10x0x0x110x0x0x1 : cnt0=17'h400;
        16'b0x10x0x110x0x0x1 : cnt0=17'h400;
        16'b1110x0x110x0x0x1 : cnt0=17'h800;
        16'b0x0x10x110x0x0x1 : cnt0=17'h400;
        16'b110x10x110x0x0x1 : cnt0=17'h800;
        16'b10x110x110x0x0x1 : cnt0=17'h800;
        16'b0x1110x110x0x0x1 : cnt0=17'h800;
        16'b111110x110x0x0x1 : cnt0=17'h1000;
        16'b0x0x0x1110x0x0x1 : cnt0=17'h400;
        16'b110x0x1110x0x0x1 : cnt0=17'h800;
        16'b10x10x1110x0x0x1 : cnt0=17'h800;
        16'b0x110x1110x0x0x1 : cnt0=17'h800;
        16'b11110x1110x0x0x1 : cnt0=17'h1000;
        16'b10x0x11110x0x0x1 : cnt0=17'h800;
        16'b0x10x11110x0x0x1 : cnt0=17'h800;
        16'b1110x11110x0x0x1 : cnt0=17'h1000;
        16'b0x0x111110x0x0x1 : cnt0=17'h800;
        16'b110x111110x0x0x1 : cnt0=17'h1000;
        16'b10x1111110x0x0x1 : cnt0=17'h1000;
        16'b0x11111110x0x0x1 : cnt0=17'h1000;
        16'b1111111110x0x0x1 : cnt0=17'h2000;
        16'b0x0x0x0x0x10x0x1 : cnt0=17'h200;
        16'b110x0x0x0x10x0x1 : cnt0=17'h400;
        16'b10x10x0x0x10x0x1 : cnt0=17'h400;
        16'b0x110x0x0x10x0x1 : cnt0=17'h400;
        16'b11110x0x0x10x0x1 : cnt0=17'h800;
        16'b10x0x10x0x10x0x1 : cnt0=17'h400;
        16'b0x10x10x0x10x0x1 : cnt0=17'h400;
        16'b1110x10x0x10x0x1 : cnt0=17'h800;
        16'b0x0x110x0x10x0x1 : cnt0=17'h400;
        16'b110x110x0x10x0x1 : cnt0=17'h800;
        16'b10x1110x0x10x0x1 : cnt0=17'h800;
        16'b0x11110x0x10x0x1 : cnt0=17'h800;
        16'b1111110x0x10x0x1 : cnt0=17'h1000;
        16'b10x0x0x10x10x0x1 : cnt0=17'h400;
        16'b0x10x0x10x10x0x1 : cnt0=17'h400;
        16'b1110x0x10x10x0x1 : cnt0=17'h800;
        16'b0x0x10x10x10x0x1 : cnt0=17'h400;
        16'b110x10x10x10x0x1 : cnt0=17'h800;
        16'b10x110x10x10x0x1 : cnt0=17'h800;
        16'b0x1110x10x10x0x1 : cnt0=17'h800;
        16'b111110x10x10x0x1 : cnt0=17'h1000;
        16'b0x0x0x110x10x0x1 : cnt0=17'h400;
        16'b110x0x110x10x0x1 : cnt0=17'h800;
        16'b10x10x110x10x0x1 : cnt0=17'h800;
        16'b0x110x110x10x0x1 : cnt0=17'h800;
        16'b11110x110x10x0x1 : cnt0=17'h1000;
        16'b10x0x1110x10x0x1 : cnt0=17'h800;
        16'b0x10x1110x10x0x1 : cnt0=17'h800;
        16'b1110x1110x10x0x1 : cnt0=17'h1000;
        16'b0x0x11110x10x0x1 : cnt0=17'h800;
        16'b110x11110x10x0x1 : cnt0=17'h1000;
        16'b10x111110x10x0x1 : cnt0=17'h1000;
        16'b0x1111110x10x0x1 : cnt0=17'h1000;
        16'b111111110x10x0x1 : cnt0=17'h2000;
        16'b10x0x0x0x110x0x1 : cnt0=17'h400;
        16'b0x10x0x0x110x0x1 : cnt0=17'h400;
        16'b1110x0x0x110x0x1 : cnt0=17'h800;
        16'b0x0x10x0x110x0x1 : cnt0=17'h400;
        16'b110x10x0x110x0x1 : cnt0=17'h800;
        16'b10x110x0x110x0x1 : cnt0=17'h800;
        16'b0x1110x0x110x0x1 : cnt0=17'h800;
        16'b111110x0x110x0x1 : cnt0=17'h1000;
        16'b0x0x0x10x110x0x1 : cnt0=17'h400;
        16'b110x0x10x110x0x1 : cnt0=17'h800;
        16'b10x10x10x110x0x1 : cnt0=17'h800;
        16'b0x110x10x110x0x1 : cnt0=17'h800;
        16'b11110x10x110x0x1 : cnt0=17'h1000;
        16'b10x0x110x110x0x1 : cnt0=17'h800;
        16'b0x10x110x110x0x1 : cnt0=17'h800;
        16'b1110x110x110x0x1 : cnt0=17'h1000;
        16'b0x0x1110x110x0x1 : cnt0=17'h800;
        16'b110x1110x110x0x1 : cnt0=17'h1000;
        16'b10x11110x110x0x1 : cnt0=17'h1000;
        16'b0x111110x110x0x1 : cnt0=17'h1000;
        16'b11111110x110x0x1 : cnt0=17'h2000;
        16'b0x0x0x0x1110x0x1 : cnt0=17'h400;
        16'b110x0x0x1110x0x1 : cnt0=17'h800;
        16'b10x10x0x1110x0x1 : cnt0=17'h800;
        16'b0x110x0x1110x0x1 : cnt0=17'h800;
        16'b11110x0x1110x0x1 : cnt0=17'h1000;
        16'b10x0x10x1110x0x1 : cnt0=17'h800;
        16'b0x10x10x1110x0x1 : cnt0=17'h800;
        16'b1110x10x1110x0x1 : cnt0=17'h1000;
        16'b0x0x110x1110x0x1 : cnt0=17'h800;
        16'b110x110x1110x0x1 : cnt0=17'h1000;
        16'b10x1110x1110x0x1 : cnt0=17'h1000;
        16'b0x11110x1110x0x1 : cnt0=17'h1000;
        16'b1111110x1110x0x1 : cnt0=17'h2000;
        16'b10x0x0x11110x0x1 : cnt0=17'h800;
        16'b0x10x0x11110x0x1 : cnt0=17'h800;
        16'b1110x0x11110x0x1 : cnt0=17'h1000;
        16'b0x0x10x11110x0x1 : cnt0=17'h800;
        16'b110x10x11110x0x1 : cnt0=17'h1000;
        16'b10x110x11110x0x1 : cnt0=17'h1000;
        16'b0x1110x11110x0x1 : cnt0=17'h1000;
        16'b111110x11110x0x1 : cnt0=17'h2000;
        16'b0x0x0x111110x0x1 : cnt0=17'h800;
        16'b110x0x111110x0x1 : cnt0=17'h1000;
        16'b10x10x111110x0x1 : cnt0=17'h1000;
        16'b0x110x111110x0x1 : cnt0=17'h1000;
        16'b11110x111110x0x1 : cnt0=17'h2000;
        16'b10x0x1111110x0x1 : cnt0=17'h1000;
        16'b0x10x1111110x0x1 : cnt0=17'h1000;
        16'b1110x1111110x0x1 : cnt0=17'h2000;
        16'b0x0x11111110x0x1 : cnt0=17'h1000;
        16'b110x11111110x0x1 : cnt0=17'h2000;
        16'b10x111111110x0x1 : cnt0=17'h2000;
        16'b0x1111111110x0x1 : cnt0=17'h2000;
        16'b111111111110x0x1 : cnt0=17'h4000;
        16'b0x0x0x0x0x0x10x1 : cnt0=17'h200;
        16'b110x0x0x0x0x10x1 : cnt0=17'h400;
        16'b10x10x0x0x0x10x1 : cnt0=17'h400;
        16'b0x110x0x0x0x10x1 : cnt0=17'h400;
        16'b11110x0x0x0x10x1 : cnt0=17'h800;
        16'b10x0x10x0x0x10x1 : cnt0=17'h400;
        16'b0x10x10x0x0x10x1 : cnt0=17'h400;
        16'b1110x10x0x0x10x1 : cnt0=17'h800;
        16'b0x0x110x0x0x10x1 : cnt0=17'h400;
        16'b110x110x0x0x10x1 : cnt0=17'h800;
        16'b10x1110x0x0x10x1 : cnt0=17'h800;
        16'b0x11110x0x0x10x1 : cnt0=17'h800;
        16'b1111110x0x0x10x1 : cnt0=17'h1000;
        16'b10x0x0x10x0x10x1 : cnt0=17'h400;
        16'b0x10x0x10x0x10x1 : cnt0=17'h400;
        16'b1110x0x10x0x10x1 : cnt0=17'h800;
        16'b0x0x10x10x0x10x1 : cnt0=17'h400;
        16'b110x10x10x0x10x1 : cnt0=17'h800;
        16'b10x110x10x0x10x1 : cnt0=17'h800;
        16'b0x1110x10x0x10x1 : cnt0=17'h800;
        16'b111110x10x0x10x1 : cnt0=17'h1000;
        16'b0x0x0x110x0x10x1 : cnt0=17'h400;
        16'b110x0x110x0x10x1 : cnt0=17'h800;
        16'b10x10x110x0x10x1 : cnt0=17'h800;
        16'b0x110x110x0x10x1 : cnt0=17'h800;
        16'b11110x110x0x10x1 : cnt0=17'h1000;
        16'b10x0x1110x0x10x1 : cnt0=17'h800;
        16'b0x10x1110x0x10x1 : cnt0=17'h800;
        16'b1110x1110x0x10x1 : cnt0=17'h1000;
        16'b0x0x11110x0x10x1 : cnt0=17'h800;
        16'b110x11110x0x10x1 : cnt0=17'h1000;
        16'b10x111110x0x10x1 : cnt0=17'h1000;
        16'b0x1111110x0x10x1 : cnt0=17'h1000;
        16'b111111110x0x10x1 : cnt0=17'h2000;
        16'b10x0x0x0x10x10x1 : cnt0=17'h400;
        16'b0x10x0x0x10x10x1 : cnt0=17'h400;
        16'b1110x0x0x10x10x1 : cnt0=17'h800;
        16'b0x0x10x0x10x10x1 : cnt0=17'h400;
        16'b110x10x0x10x10x1 : cnt0=17'h800;
        16'b10x110x0x10x10x1 : cnt0=17'h800;
        16'b0x1110x0x10x10x1 : cnt0=17'h800;
        16'b111110x0x10x10x1 : cnt0=17'h1000;
        16'b0x0x0x10x10x10x1 : cnt0=17'h400;
        16'b110x0x10x10x10x1 : cnt0=17'h800;
        16'b10x10x10x10x10x1 : cnt0=17'h800;
        16'b0x110x10x10x10x1 : cnt0=17'h800;
        16'b11110x10x10x10x1 : cnt0=17'h1000;
        16'b10x0x110x10x10x1 : cnt0=17'h800;
        16'b0x10x110x10x10x1 : cnt0=17'h800;
        16'b1110x110x10x10x1 : cnt0=17'h1000;
        16'b0x0x1110x10x10x1 : cnt0=17'h800;
        16'b110x1110x10x10x1 : cnt0=17'h1000;
        16'b10x11110x10x10x1 : cnt0=17'h1000;
        16'b0x111110x10x10x1 : cnt0=17'h1000;
        16'b11111110x10x10x1 : cnt0=17'h2000;
        16'b0x0x0x0x110x10x1 : cnt0=17'h400;
        16'b110x0x0x110x10x1 : cnt0=17'h800;
        16'b10x10x0x110x10x1 : cnt0=17'h800;
        16'b0x110x0x110x10x1 : cnt0=17'h800;
        16'b11110x0x110x10x1 : cnt0=17'h1000;
        16'b10x0x10x110x10x1 : cnt0=17'h800;
        16'b0x10x10x110x10x1 : cnt0=17'h800;
        16'b1110x10x110x10x1 : cnt0=17'h1000;
        16'b0x0x110x110x10x1 : cnt0=17'h800;
        16'b110x110x110x10x1 : cnt0=17'h1000;
        16'b10x1110x110x10x1 : cnt0=17'h1000;
        16'b0x11110x110x10x1 : cnt0=17'h1000;
        16'b1111110x110x10x1 : cnt0=17'h2000;
        16'b10x0x0x1110x10x1 : cnt0=17'h800;
        16'b0x10x0x1110x10x1 : cnt0=17'h800;
        16'b1110x0x1110x10x1 : cnt0=17'h1000;
        16'b0x0x10x1110x10x1 : cnt0=17'h800;
        16'b110x10x1110x10x1 : cnt0=17'h1000;
        16'b10x110x1110x10x1 : cnt0=17'h1000;
        16'b0x1110x1110x10x1 : cnt0=17'h1000;
        16'b111110x1110x10x1 : cnt0=17'h2000;
        16'b0x0x0x11110x10x1 : cnt0=17'h800;
        16'b110x0x11110x10x1 : cnt0=17'h1000;
        16'b10x10x11110x10x1 : cnt0=17'h1000;
        16'b0x110x11110x10x1 : cnt0=17'h1000;
        16'b11110x11110x10x1 : cnt0=17'h2000;
        16'b10x0x111110x10x1 : cnt0=17'h1000;
        16'b0x10x111110x10x1 : cnt0=17'h1000;
        16'b1110x111110x10x1 : cnt0=17'h2000;
        16'b0x0x1111110x10x1 : cnt0=17'h1000;
        16'b110x1111110x10x1 : cnt0=17'h2000;
        16'b10x11111110x10x1 : cnt0=17'h2000;
        16'b0x111111110x10x1 : cnt0=17'h2000;
        16'b11111111110x10x1 : cnt0=17'h4000;
        16'b10x0x0x0x0x110x1 : cnt0=17'h400;
        16'b0x10x0x0x0x110x1 : cnt0=17'h400;
        16'b1110x0x0x0x110x1 : cnt0=17'h800;
        16'b0x0x10x0x0x110x1 : cnt0=17'h400;
        16'b110x10x0x0x110x1 : cnt0=17'h800;
        16'b10x110x0x0x110x1 : cnt0=17'h800;
        16'b0x1110x0x0x110x1 : cnt0=17'h800;
        16'b111110x0x0x110x1 : cnt0=17'h1000;
        16'b0x0x0x10x0x110x1 : cnt0=17'h400;
        16'b110x0x10x0x110x1 : cnt0=17'h800;
        16'b10x10x10x0x110x1 : cnt0=17'h800;
        16'b0x110x10x0x110x1 : cnt0=17'h800;
        16'b11110x10x0x110x1 : cnt0=17'h1000;
        16'b10x0x110x0x110x1 : cnt0=17'h800;
        16'b0x10x110x0x110x1 : cnt0=17'h800;
        16'b1110x110x0x110x1 : cnt0=17'h1000;
        16'b0x0x1110x0x110x1 : cnt0=17'h800;
        16'b110x1110x0x110x1 : cnt0=17'h1000;
        16'b10x11110x0x110x1 : cnt0=17'h1000;
        16'b0x111110x0x110x1 : cnt0=17'h1000;
        16'b11111110x0x110x1 : cnt0=17'h2000;
        16'b0x0x0x0x10x110x1 : cnt0=17'h400;
        16'b110x0x0x10x110x1 : cnt0=17'h800;
        16'b10x10x0x10x110x1 : cnt0=17'h800;
        16'b0x110x0x10x110x1 : cnt0=17'h800;
        16'b11110x0x10x110x1 : cnt0=17'h1000;
        16'b10x0x10x10x110x1 : cnt0=17'h800;
        16'b0x10x10x10x110x1 : cnt0=17'h800;
        16'b1110x10x10x110x1 : cnt0=17'h1000;
        16'b0x0x110x10x110x1 : cnt0=17'h800;
        16'b110x110x10x110x1 : cnt0=17'h1000;
        16'b10x1110x10x110x1 : cnt0=17'h1000;
        16'b0x11110x10x110x1 : cnt0=17'h1000;
        16'b1111110x10x110x1 : cnt0=17'h2000;
        16'b10x0x0x110x110x1 : cnt0=17'h800;
        16'b0x10x0x110x110x1 : cnt0=17'h800;
        16'b1110x0x110x110x1 : cnt0=17'h1000;
        16'b0x0x10x110x110x1 : cnt0=17'h800;
        16'b110x10x110x110x1 : cnt0=17'h1000;
        16'b10x110x110x110x1 : cnt0=17'h1000;
        16'b0x1110x110x110x1 : cnt0=17'h1000;
        16'b111110x110x110x1 : cnt0=17'h2000;
        16'b0x0x0x1110x110x1 : cnt0=17'h800;
        16'b110x0x1110x110x1 : cnt0=17'h1000;
        16'b10x10x1110x110x1 : cnt0=17'h1000;
        16'b0x110x1110x110x1 : cnt0=17'h1000;
        16'b11110x1110x110x1 : cnt0=17'h2000;
        16'b10x0x11110x110x1 : cnt0=17'h1000;
        16'b0x10x11110x110x1 : cnt0=17'h1000;
        16'b1110x11110x110x1 : cnt0=17'h2000;
        16'b0x0x111110x110x1 : cnt0=17'h1000;
        16'b110x111110x110x1 : cnt0=17'h2000;
        16'b10x1111110x110x1 : cnt0=17'h2000;
        16'b0x11111110x110x1 : cnt0=17'h2000;
        16'b1111111110x110x1 : cnt0=17'h4000;
        16'b0x0x0x0x0x1110x1 : cnt0=17'h400;
        16'b110x0x0x0x1110x1 : cnt0=17'h800;
        16'b10x10x0x0x1110x1 : cnt0=17'h800;
        16'b0x110x0x0x1110x1 : cnt0=17'h800;
        16'b11110x0x0x1110x1 : cnt0=17'h1000;
        16'b10x0x10x0x1110x1 : cnt0=17'h800;
        16'b0x10x10x0x1110x1 : cnt0=17'h800;
        16'b1110x10x0x1110x1 : cnt0=17'h1000;
        16'b0x0x110x0x1110x1 : cnt0=17'h800;
        16'b110x110x0x1110x1 : cnt0=17'h1000;
        16'b10x1110x0x1110x1 : cnt0=17'h1000;
        16'b0x11110x0x1110x1 : cnt0=17'h1000;
        16'b1111110x0x1110x1 : cnt0=17'h2000;
        16'b10x0x0x10x1110x1 : cnt0=17'h800;
        16'b0x10x0x10x1110x1 : cnt0=17'h800;
        16'b1110x0x10x1110x1 : cnt0=17'h1000;
        16'b0x0x10x10x1110x1 : cnt0=17'h800;
        16'b110x10x10x1110x1 : cnt0=17'h1000;
        16'b10x110x10x1110x1 : cnt0=17'h1000;
        16'b0x1110x10x1110x1 : cnt0=17'h1000;
        16'b111110x10x1110x1 : cnt0=17'h2000;
        16'b0x0x0x110x1110x1 : cnt0=17'h800;
        16'b110x0x110x1110x1 : cnt0=17'h1000;
        16'b10x10x110x1110x1 : cnt0=17'h1000;
        16'b0x110x110x1110x1 : cnt0=17'h1000;
        16'b11110x110x1110x1 : cnt0=17'h2000;
        16'b10x0x1110x1110x1 : cnt0=17'h1000;
        16'b0x10x1110x1110x1 : cnt0=17'h1000;
        16'b1110x1110x1110x1 : cnt0=17'h2000;
        16'b0x0x11110x1110x1 : cnt0=17'h1000;
        16'b110x11110x1110x1 : cnt0=17'h2000;
        16'b10x111110x1110x1 : cnt0=17'h2000;
        16'b0x1111110x1110x1 : cnt0=17'h2000;
        16'b111111110x1110x1 : cnt0=17'h4000;
        16'b10x0x0x0x11110x1 : cnt0=17'h800;
        16'b0x10x0x0x11110x1 : cnt0=17'h800;
        16'b1110x0x0x11110x1 : cnt0=17'h1000;
        16'b0x0x10x0x11110x1 : cnt0=17'h800;
        16'b110x10x0x11110x1 : cnt0=17'h1000;
        16'b10x110x0x11110x1 : cnt0=17'h1000;
        16'b0x1110x0x11110x1 : cnt0=17'h1000;
        16'b111110x0x11110x1 : cnt0=17'h2000;
        16'b0x0x0x10x11110x1 : cnt0=17'h800;
        16'b110x0x10x11110x1 : cnt0=17'h1000;
        16'b10x10x10x11110x1 : cnt0=17'h1000;
        16'b0x110x10x11110x1 : cnt0=17'h1000;
        16'b11110x10x11110x1 : cnt0=17'h2000;
        16'b10x0x110x11110x1 : cnt0=17'h1000;
        16'b0x10x110x11110x1 : cnt0=17'h1000;
        16'b1110x110x11110x1 : cnt0=17'h2000;
        16'b0x0x1110x11110x1 : cnt0=17'h1000;
        16'b110x1110x11110x1 : cnt0=17'h2000;
        16'b10x11110x11110x1 : cnt0=17'h2000;
        16'b0x111110x11110x1 : cnt0=17'h2000;
        16'b11111110x11110x1 : cnt0=17'h4000;
        16'b0x0x0x0x111110x1 : cnt0=17'h800;
        16'b110x0x0x111110x1 : cnt0=17'h1000;
        16'b10x10x0x111110x1 : cnt0=17'h1000;
        16'b0x110x0x111110x1 : cnt0=17'h1000;
        16'b11110x0x111110x1 : cnt0=17'h2000;
        16'b10x0x10x111110x1 : cnt0=17'h1000;
        16'b0x10x10x111110x1 : cnt0=17'h1000;
        16'b1110x10x111110x1 : cnt0=17'h2000;
        16'b0x0x110x111110x1 : cnt0=17'h1000;
        16'b110x110x111110x1 : cnt0=17'h2000;
        16'b10x1110x111110x1 : cnt0=17'h2000;
        16'b0x11110x111110x1 : cnt0=17'h2000;
        16'b1111110x111110x1 : cnt0=17'h4000;
        16'b10x0x0x1111110x1 : cnt0=17'h1000;
        16'b0x10x0x1111110x1 : cnt0=17'h1000;
        16'b1110x0x1111110x1 : cnt0=17'h2000;
        16'b0x0x10x1111110x1 : cnt0=17'h1000;
        16'b110x10x1111110x1 : cnt0=17'h2000;
        16'b10x110x1111110x1 : cnt0=17'h2000;
        16'b0x1110x1111110x1 : cnt0=17'h2000;
        16'b111110x1111110x1 : cnt0=17'h4000;
        16'b0x0x0x11111110x1 : cnt0=17'h1000;
        16'b110x0x11111110x1 : cnt0=17'h2000;
        16'b10x10x11111110x1 : cnt0=17'h2000;
        16'b0x110x11111110x1 : cnt0=17'h2000;
        16'b11110x11111110x1 : cnt0=17'h4000;
        16'b10x0x111111110x1 : cnt0=17'h2000;
        16'b0x10x111111110x1 : cnt0=17'h2000;
        16'b1110x111111110x1 : cnt0=17'h4000;
        16'b0x0x1111111110x1 : cnt0=17'h2000;
        16'b110x1111111110x1 : cnt0=17'h4000;
        16'b10x11111111110x1 : cnt0=17'h4000;
        16'b0x111111111110x1 : cnt0=17'h4000;
        16'b11111111111110x1 : cnt0=17'h8000;
        16'b0x0x0x0x0x0x0x11 : cnt0=17'h200;
        16'b110x0x0x0x0x0x11 : cnt0=17'h400;
        16'b10x10x0x0x0x0x11 : cnt0=17'h400;
        16'b0x110x0x0x0x0x11 : cnt0=17'h400;
        16'b11110x0x0x0x0x11 : cnt0=17'h800;
        16'b10x0x10x0x0x0x11 : cnt0=17'h400;
        16'b0x10x10x0x0x0x11 : cnt0=17'h400;
        16'b1110x10x0x0x0x11 : cnt0=17'h800;
        16'b0x0x110x0x0x0x11 : cnt0=17'h400;
        16'b110x110x0x0x0x11 : cnt0=17'h800;
        16'b10x1110x0x0x0x11 : cnt0=17'h800;
        16'b0x11110x0x0x0x11 : cnt0=17'h800;
        16'b1111110x0x0x0x11 : cnt0=17'h1000;
        16'b10x0x0x10x0x0x11 : cnt0=17'h400;
        16'b0x10x0x10x0x0x11 : cnt0=17'h400;
        16'b1110x0x10x0x0x11 : cnt0=17'h800;
        16'b0x0x10x10x0x0x11 : cnt0=17'h400;
        16'b110x10x10x0x0x11 : cnt0=17'h800;
        16'b10x110x10x0x0x11 : cnt0=17'h800;
        16'b0x1110x10x0x0x11 : cnt0=17'h800;
        16'b111110x10x0x0x11 : cnt0=17'h1000;
        16'b0x0x0x110x0x0x11 : cnt0=17'h400;
        16'b110x0x110x0x0x11 : cnt0=17'h800;
        16'b10x10x110x0x0x11 : cnt0=17'h800;
        16'b0x110x110x0x0x11 : cnt0=17'h800;
        16'b11110x110x0x0x11 : cnt0=17'h1000;
        16'b10x0x1110x0x0x11 : cnt0=17'h800;
        16'b0x10x1110x0x0x11 : cnt0=17'h800;
        16'b1110x1110x0x0x11 : cnt0=17'h1000;
        16'b0x0x11110x0x0x11 : cnt0=17'h800;
        16'b110x11110x0x0x11 : cnt0=17'h1000;
        16'b10x111110x0x0x11 : cnt0=17'h1000;
        16'b0x1111110x0x0x11 : cnt0=17'h1000;
        16'b111111110x0x0x11 : cnt0=17'h2000;
        16'b10x0x0x0x10x0x11 : cnt0=17'h400;
        16'b0x10x0x0x10x0x11 : cnt0=17'h400;
        16'b1110x0x0x10x0x11 : cnt0=17'h800;
        16'b0x0x10x0x10x0x11 : cnt0=17'h400;
        16'b110x10x0x10x0x11 : cnt0=17'h800;
        16'b10x110x0x10x0x11 : cnt0=17'h800;
        16'b0x1110x0x10x0x11 : cnt0=17'h800;
        16'b111110x0x10x0x11 : cnt0=17'h1000;
        16'b0x0x0x10x10x0x11 : cnt0=17'h400;
        16'b110x0x10x10x0x11 : cnt0=17'h800;
        16'b10x10x10x10x0x11 : cnt0=17'h800;
        16'b0x110x10x10x0x11 : cnt0=17'h800;
        16'b11110x10x10x0x11 : cnt0=17'h1000;
        16'b10x0x110x10x0x11 : cnt0=17'h800;
        16'b0x10x110x10x0x11 : cnt0=17'h800;
        16'b1110x110x10x0x11 : cnt0=17'h1000;
        16'b0x0x1110x10x0x11 : cnt0=17'h800;
        16'b110x1110x10x0x11 : cnt0=17'h1000;
        16'b10x11110x10x0x11 : cnt0=17'h1000;
        16'b0x111110x10x0x11 : cnt0=17'h1000;
        16'b11111110x10x0x11 : cnt0=17'h2000;
        16'b0x0x0x0x110x0x11 : cnt0=17'h400;
        16'b110x0x0x110x0x11 : cnt0=17'h800;
        16'b10x10x0x110x0x11 : cnt0=17'h800;
        16'b0x110x0x110x0x11 : cnt0=17'h800;
        16'b11110x0x110x0x11 : cnt0=17'h1000;
        16'b10x0x10x110x0x11 : cnt0=17'h800;
        16'b0x10x10x110x0x11 : cnt0=17'h800;
        16'b1110x10x110x0x11 : cnt0=17'h1000;
        16'b0x0x110x110x0x11 : cnt0=17'h800;
        16'b110x110x110x0x11 : cnt0=17'h1000;
        16'b10x1110x110x0x11 : cnt0=17'h1000;
        16'b0x11110x110x0x11 : cnt0=17'h1000;
        16'b1111110x110x0x11 : cnt0=17'h2000;
        16'b10x0x0x1110x0x11 : cnt0=17'h800;
        16'b0x10x0x1110x0x11 : cnt0=17'h800;
        16'b1110x0x1110x0x11 : cnt0=17'h1000;
        16'b0x0x10x1110x0x11 : cnt0=17'h800;
        16'b110x10x1110x0x11 : cnt0=17'h1000;
        16'b10x110x1110x0x11 : cnt0=17'h1000;
        16'b0x1110x1110x0x11 : cnt0=17'h1000;
        16'b111110x1110x0x11 : cnt0=17'h2000;
        16'b0x0x0x11110x0x11 : cnt0=17'h800;
        16'b110x0x11110x0x11 : cnt0=17'h1000;
        16'b10x10x11110x0x11 : cnt0=17'h1000;
        16'b0x110x11110x0x11 : cnt0=17'h1000;
        16'b11110x11110x0x11 : cnt0=17'h2000;
        16'b10x0x111110x0x11 : cnt0=17'h1000;
        16'b0x10x111110x0x11 : cnt0=17'h1000;
        16'b1110x111110x0x11 : cnt0=17'h2000;
        16'b0x0x1111110x0x11 : cnt0=17'h1000;
        16'b110x1111110x0x11 : cnt0=17'h2000;
        16'b10x11111110x0x11 : cnt0=17'h2000;
        16'b0x111111110x0x11 : cnt0=17'h2000;
        16'b11111111110x0x11 : cnt0=17'h4000;
        16'b10x0x0x0x0x10x11 : cnt0=17'h400;
        16'b0x10x0x0x0x10x11 : cnt0=17'h400;
        16'b1110x0x0x0x10x11 : cnt0=17'h800;
        16'b0x0x10x0x0x10x11 : cnt0=17'h400;
        16'b110x10x0x0x10x11 : cnt0=17'h800;
        16'b10x110x0x0x10x11 : cnt0=17'h800;
        16'b0x1110x0x0x10x11 : cnt0=17'h800;
        16'b111110x0x0x10x11 : cnt0=17'h1000;
        16'b0x0x0x10x0x10x11 : cnt0=17'h400;
        16'b110x0x10x0x10x11 : cnt0=17'h800;
        16'b10x10x10x0x10x11 : cnt0=17'h800;
        16'b0x110x10x0x10x11 : cnt0=17'h800;
        16'b11110x10x0x10x11 : cnt0=17'h1000;
        16'b10x0x110x0x10x11 : cnt0=17'h800;
        16'b0x10x110x0x10x11 : cnt0=17'h800;
        16'b1110x110x0x10x11 : cnt0=17'h1000;
        16'b0x0x1110x0x10x11 : cnt0=17'h800;
        16'b110x1110x0x10x11 : cnt0=17'h1000;
        16'b10x11110x0x10x11 : cnt0=17'h1000;
        16'b0x111110x0x10x11 : cnt0=17'h1000;
        16'b11111110x0x10x11 : cnt0=17'h2000;
        16'b0x0x0x0x10x10x11 : cnt0=17'h400;
        16'b110x0x0x10x10x11 : cnt0=17'h800;
        16'b10x10x0x10x10x11 : cnt0=17'h800;
        16'b0x110x0x10x10x11 : cnt0=17'h800;
        16'b11110x0x10x10x11 : cnt0=17'h1000;
        16'b10x0x10x10x10x11 : cnt0=17'h800;
        16'b0x10x10x10x10x11 : cnt0=17'h800;
        16'b1110x10x10x10x11 : cnt0=17'h1000;
        16'b0x0x110x10x10x11 : cnt0=17'h800;
        16'b110x110x10x10x11 : cnt0=17'h1000;
        16'b10x1110x10x10x11 : cnt0=17'h1000;
        16'b0x11110x10x10x11 : cnt0=17'h1000;
        16'b1111110x10x10x11 : cnt0=17'h2000;
        16'b10x0x0x110x10x11 : cnt0=17'h800;
        16'b0x10x0x110x10x11 : cnt0=17'h800;
        16'b1110x0x110x10x11 : cnt0=17'h1000;
        16'b0x0x10x110x10x11 : cnt0=17'h800;
        16'b110x10x110x10x11 : cnt0=17'h1000;
        16'b10x110x110x10x11 : cnt0=17'h1000;
        16'b0x1110x110x10x11 : cnt0=17'h1000;
        16'b111110x110x10x11 : cnt0=17'h2000;
        16'b0x0x0x1110x10x11 : cnt0=17'h800;
        16'b110x0x1110x10x11 : cnt0=17'h1000;
        16'b10x10x1110x10x11 : cnt0=17'h1000;
        16'b0x110x1110x10x11 : cnt0=17'h1000;
        16'b11110x1110x10x11 : cnt0=17'h2000;
        16'b10x0x11110x10x11 : cnt0=17'h1000;
        16'b0x10x11110x10x11 : cnt0=17'h1000;
        16'b1110x11110x10x11 : cnt0=17'h2000;
        16'b0x0x111110x10x11 : cnt0=17'h1000;
        16'b110x111110x10x11 : cnt0=17'h2000;
        16'b10x1111110x10x11 : cnt0=17'h2000;
        16'b0x11111110x10x11 : cnt0=17'h2000;
        16'b1111111110x10x11 : cnt0=17'h4000;
        16'b0x0x0x0x0x110x11 : cnt0=17'h400;
        16'b110x0x0x0x110x11 : cnt0=17'h800;
        16'b10x10x0x0x110x11 : cnt0=17'h800;
        16'b0x110x0x0x110x11 : cnt0=17'h800;
        16'b11110x0x0x110x11 : cnt0=17'h1000;
        16'b10x0x10x0x110x11 : cnt0=17'h800;
        16'b0x10x10x0x110x11 : cnt0=17'h800;
        16'b1110x10x0x110x11 : cnt0=17'h1000;
        16'b0x0x110x0x110x11 : cnt0=17'h800;
        16'b110x110x0x110x11 : cnt0=17'h1000;
        16'b10x1110x0x110x11 : cnt0=17'h1000;
        16'b0x11110x0x110x11 : cnt0=17'h1000;
        16'b1111110x0x110x11 : cnt0=17'h2000;
        16'b10x0x0x10x110x11 : cnt0=17'h800;
        16'b0x10x0x10x110x11 : cnt0=17'h800;
        16'b1110x0x10x110x11 : cnt0=17'h1000;
        16'b0x0x10x10x110x11 : cnt0=17'h800;
        16'b110x10x10x110x11 : cnt0=17'h1000;
        16'b10x110x10x110x11 : cnt0=17'h1000;
        16'b0x1110x10x110x11 : cnt0=17'h1000;
        16'b111110x10x110x11 : cnt0=17'h2000;
        16'b0x0x0x110x110x11 : cnt0=17'h800;
        16'b110x0x110x110x11 : cnt0=17'h1000;
        16'b10x10x110x110x11 : cnt0=17'h1000;
        16'b0x110x110x110x11 : cnt0=17'h1000;
        16'b11110x110x110x11 : cnt0=17'h2000;
        16'b10x0x1110x110x11 : cnt0=17'h1000;
        16'b0x10x1110x110x11 : cnt0=17'h1000;
        16'b1110x1110x110x11 : cnt0=17'h2000;
        16'b0x0x11110x110x11 : cnt0=17'h1000;
        16'b110x11110x110x11 : cnt0=17'h2000;
        16'b10x111110x110x11 : cnt0=17'h2000;
        16'b0x1111110x110x11 : cnt0=17'h2000;
        16'b111111110x110x11 : cnt0=17'h4000;
        16'b10x0x0x0x1110x11 : cnt0=17'h800;
        16'b0x10x0x0x1110x11 : cnt0=17'h800;
        16'b1110x0x0x1110x11 : cnt0=17'h1000;
        16'b0x0x10x0x1110x11 : cnt0=17'h800;
        16'b110x10x0x1110x11 : cnt0=17'h1000;
        16'b10x110x0x1110x11 : cnt0=17'h1000;
        16'b0x1110x0x1110x11 : cnt0=17'h1000;
        16'b111110x0x1110x11 : cnt0=17'h2000;
        16'b0x0x0x10x1110x11 : cnt0=17'h800;
        16'b110x0x10x1110x11 : cnt0=17'h1000;
        16'b10x10x10x1110x11 : cnt0=17'h1000;
        16'b0x110x10x1110x11 : cnt0=17'h1000;
        16'b11110x10x1110x11 : cnt0=17'h2000;
        16'b10x0x110x1110x11 : cnt0=17'h1000;
        16'b0x10x110x1110x11 : cnt0=17'h1000;
        16'b1110x110x1110x11 : cnt0=17'h2000;
        16'b0x0x1110x1110x11 : cnt0=17'h1000;
        16'b110x1110x1110x11 : cnt0=17'h2000;
        16'b10x11110x1110x11 : cnt0=17'h2000;
        16'b0x111110x1110x11 : cnt0=17'h2000;
        16'b11111110x1110x11 : cnt0=17'h4000;
        16'b0x0x0x0x11110x11 : cnt0=17'h800;
        16'b110x0x0x11110x11 : cnt0=17'h1000;
        16'b10x10x0x11110x11 : cnt0=17'h1000;
        16'b0x110x0x11110x11 : cnt0=17'h1000;
        16'b11110x0x11110x11 : cnt0=17'h2000;
        16'b10x0x10x11110x11 : cnt0=17'h1000;
        16'b0x10x10x11110x11 : cnt0=17'h1000;
        16'b1110x10x11110x11 : cnt0=17'h2000;
        16'b0x0x110x11110x11 : cnt0=17'h1000;
        16'b110x110x11110x11 : cnt0=17'h2000;
        16'b10x1110x11110x11 : cnt0=17'h2000;
        16'b0x11110x11110x11 : cnt0=17'h2000;
        16'b1111110x11110x11 : cnt0=17'h4000;
        16'b10x0x0x111110x11 : cnt0=17'h1000;
        16'b0x10x0x111110x11 : cnt0=17'h1000;
        16'b1110x0x111110x11 : cnt0=17'h2000;
        16'b0x0x10x111110x11 : cnt0=17'h1000;
        16'b110x10x111110x11 : cnt0=17'h2000;
        16'b10x110x111110x11 : cnt0=17'h2000;
        16'b0x1110x111110x11 : cnt0=17'h2000;
        16'b111110x111110x11 : cnt0=17'h4000;
        16'b0x0x0x1111110x11 : cnt0=17'h1000;
        16'b110x0x1111110x11 : cnt0=17'h2000;
        16'b10x10x1111110x11 : cnt0=17'h2000;
        16'b0x110x1111110x11 : cnt0=17'h2000;
        16'b11110x1111110x11 : cnt0=17'h4000;
        16'b10x0x11111110x11 : cnt0=17'h2000;
        16'b0x10x11111110x11 : cnt0=17'h2000;
        16'b1110x11111110x11 : cnt0=17'h4000;
        16'b0x0x111111110x11 : cnt0=17'h2000;
        16'b110x111111110x11 : cnt0=17'h4000;
        16'b10x1111111110x11 : cnt0=17'h4000;
        16'b0x11111111110x11 : cnt0=17'h4000;
        16'b1111111111110x11 : cnt0=17'h8000;
        16'b10x0x0x0x0x0x111 : cnt0=17'h400;
        16'b0x10x0x0x0x0x111 : cnt0=17'h400;
        16'b1110x0x0x0x0x111 : cnt0=17'h800;
        16'b0x0x10x0x0x0x111 : cnt0=17'h400;
        16'b110x10x0x0x0x111 : cnt0=17'h800;
        16'b10x110x0x0x0x111 : cnt0=17'h800;
        16'b0x1110x0x0x0x111 : cnt0=17'h800;
        16'b111110x0x0x0x111 : cnt0=17'h1000;
        16'b0x0x0x10x0x0x111 : cnt0=17'h400;
        16'b110x0x10x0x0x111 : cnt0=17'h800;
        16'b10x10x10x0x0x111 : cnt0=17'h800;
        16'b0x110x10x0x0x111 : cnt0=17'h800;
        16'b11110x10x0x0x111 : cnt0=17'h1000;
        16'b10x0x110x0x0x111 : cnt0=17'h800;
        16'b0x10x110x0x0x111 : cnt0=17'h800;
        16'b1110x110x0x0x111 : cnt0=17'h1000;
        16'b0x0x1110x0x0x111 : cnt0=17'h800;
        16'b110x1110x0x0x111 : cnt0=17'h1000;
        16'b10x11110x0x0x111 : cnt0=17'h1000;
        16'b0x111110x0x0x111 : cnt0=17'h1000;
        16'b11111110x0x0x111 : cnt0=17'h2000;
        16'b0x0x0x0x10x0x111 : cnt0=17'h400;
        16'b110x0x0x10x0x111 : cnt0=17'h800;
        16'b10x10x0x10x0x111 : cnt0=17'h800;
        16'b0x110x0x10x0x111 : cnt0=17'h800;
        16'b11110x0x10x0x111 : cnt0=17'h1000;
        16'b10x0x10x10x0x111 : cnt0=17'h800;
        16'b0x10x10x10x0x111 : cnt0=17'h800;
        16'b1110x10x10x0x111 : cnt0=17'h1000;
        16'b0x0x110x10x0x111 : cnt0=17'h800;
        16'b110x110x10x0x111 : cnt0=17'h1000;
        16'b10x1110x10x0x111 : cnt0=17'h1000;
        16'b0x11110x10x0x111 : cnt0=17'h1000;
        16'b1111110x10x0x111 : cnt0=17'h2000;
        16'b10x0x0x110x0x111 : cnt0=17'h800;
        16'b0x10x0x110x0x111 : cnt0=17'h800;
        16'b1110x0x110x0x111 : cnt0=17'h1000;
        16'b0x0x10x110x0x111 : cnt0=17'h800;
        16'b110x10x110x0x111 : cnt0=17'h1000;
        16'b10x110x110x0x111 : cnt0=17'h1000;
        16'b0x1110x110x0x111 : cnt0=17'h1000;
        16'b111110x110x0x111 : cnt0=17'h2000;
        16'b0x0x0x1110x0x111 : cnt0=17'h800;
        16'b110x0x1110x0x111 : cnt0=17'h1000;
        16'b10x10x1110x0x111 : cnt0=17'h1000;
        16'b0x110x1110x0x111 : cnt0=17'h1000;
        16'b11110x1110x0x111 : cnt0=17'h2000;
        16'b10x0x11110x0x111 : cnt0=17'h1000;
        16'b0x10x11110x0x111 : cnt0=17'h1000;
        16'b1110x11110x0x111 : cnt0=17'h2000;
        16'b0x0x111110x0x111 : cnt0=17'h1000;
        16'b110x111110x0x111 : cnt0=17'h2000;
        16'b10x1111110x0x111 : cnt0=17'h2000;
        16'b0x11111110x0x111 : cnt0=17'h2000;
        16'b1111111110x0x111 : cnt0=17'h4000;
        16'b0x0x0x0x0x10x111 : cnt0=17'h400;
        16'b110x0x0x0x10x111 : cnt0=17'h800;
        16'b10x10x0x0x10x111 : cnt0=17'h800;
        16'b0x110x0x0x10x111 : cnt0=17'h800;
        16'b11110x0x0x10x111 : cnt0=17'h1000;
        16'b10x0x10x0x10x111 : cnt0=17'h800;
        16'b0x10x10x0x10x111 : cnt0=17'h800;
        16'b1110x10x0x10x111 : cnt0=17'h1000;
        16'b0x0x110x0x10x111 : cnt0=17'h800;
        16'b110x110x0x10x111 : cnt0=17'h1000;
        16'b10x1110x0x10x111 : cnt0=17'h1000;
        16'b0x11110x0x10x111 : cnt0=17'h1000;
        16'b1111110x0x10x111 : cnt0=17'h2000;
        16'b10x0x0x10x10x111 : cnt0=17'h800;
        16'b0x10x0x10x10x111 : cnt0=17'h800;
        16'b1110x0x10x10x111 : cnt0=17'h1000;
        16'b0x0x10x10x10x111 : cnt0=17'h800;
        16'b110x10x10x10x111 : cnt0=17'h1000;
        16'b10x110x10x10x111 : cnt0=17'h1000;
        16'b0x1110x10x10x111 : cnt0=17'h1000;
        16'b111110x10x10x111 : cnt0=17'h2000;
        16'b0x0x0x110x10x111 : cnt0=17'h800;
        16'b110x0x110x10x111 : cnt0=17'h1000;
        16'b10x10x110x10x111 : cnt0=17'h1000;
        16'b0x110x110x10x111 : cnt0=17'h1000;
        16'b11110x110x10x111 : cnt0=17'h2000;
        16'b10x0x1110x10x111 : cnt0=17'h1000;
        16'b0x10x1110x10x111 : cnt0=17'h1000;
        16'b1110x1110x10x111 : cnt0=17'h2000;
        16'b0x0x11110x10x111 : cnt0=17'h1000;
        16'b110x11110x10x111 : cnt0=17'h2000;
        16'b10x111110x10x111 : cnt0=17'h2000;
        16'b0x1111110x10x111 : cnt0=17'h2000;
        16'b111111110x10x111 : cnt0=17'h4000;
        16'b10x0x0x0x110x111 : cnt0=17'h800;
        16'b0x10x0x0x110x111 : cnt0=17'h800;
        16'b1110x0x0x110x111 : cnt0=17'h1000;
        16'b0x0x10x0x110x111 : cnt0=17'h800;
        16'b110x10x0x110x111 : cnt0=17'h1000;
        16'b10x110x0x110x111 : cnt0=17'h1000;
        16'b0x1110x0x110x111 : cnt0=17'h1000;
        16'b111110x0x110x111 : cnt0=17'h2000;
        16'b0x0x0x10x110x111 : cnt0=17'h800;
        16'b110x0x10x110x111 : cnt0=17'h1000;
        16'b10x10x10x110x111 : cnt0=17'h1000;
        16'b0x110x10x110x111 : cnt0=17'h1000;
        16'b11110x10x110x111 : cnt0=17'h2000;
        16'b10x0x110x110x111 : cnt0=17'h1000;
        16'b0x10x110x110x111 : cnt0=17'h1000;
        16'b1110x110x110x111 : cnt0=17'h2000;
        16'b0x0x1110x110x111 : cnt0=17'h1000;
        16'b110x1110x110x111 : cnt0=17'h2000;
        16'b10x11110x110x111 : cnt0=17'h2000;
        16'b0x111110x110x111 : cnt0=17'h2000;
        16'b11111110x110x111 : cnt0=17'h4000;
        16'b0x0x0x0x1110x111 : cnt0=17'h800;
        16'b110x0x0x1110x111 : cnt0=17'h1000;
        16'b10x10x0x1110x111 : cnt0=17'h1000;
        16'b0x110x0x1110x111 : cnt0=17'h1000;
        16'b11110x0x1110x111 : cnt0=17'h2000;
        16'b10x0x10x1110x111 : cnt0=17'h1000;
        16'b0x10x10x1110x111 : cnt0=17'h1000;
        16'b1110x10x1110x111 : cnt0=17'h2000;
        16'b0x0x110x1110x111 : cnt0=17'h1000;
        16'b110x110x1110x111 : cnt0=17'h2000;
        16'b10x1110x1110x111 : cnt0=17'h2000;
        16'b0x11110x1110x111 : cnt0=17'h2000;
        16'b1111110x1110x111 : cnt0=17'h4000;
        16'b10x0x0x11110x111 : cnt0=17'h1000;
        16'b0x10x0x11110x111 : cnt0=17'h1000;
        16'b1110x0x11110x111 : cnt0=17'h2000;
        16'b0x0x10x11110x111 : cnt0=17'h1000;
        16'b110x10x11110x111 : cnt0=17'h2000;
        16'b10x110x11110x111 : cnt0=17'h2000;
        16'b0x1110x11110x111 : cnt0=17'h2000;
        16'b111110x11110x111 : cnt0=17'h4000;
        16'b0x0x0x111110x111 : cnt0=17'h1000;
        16'b110x0x111110x111 : cnt0=17'h2000;
        16'b10x10x111110x111 : cnt0=17'h2000;
        16'b0x110x111110x111 : cnt0=17'h2000;
        16'b11110x111110x111 : cnt0=17'h4000;
        16'b10x0x1111110x111 : cnt0=17'h2000;
        16'b0x10x1111110x111 : cnt0=17'h2000;
        16'b1110x1111110x111 : cnt0=17'h4000;
        16'b0x0x11111110x111 : cnt0=17'h2000;
        16'b110x11111110x111 : cnt0=17'h4000;
        16'b10x111111110x111 : cnt0=17'h4000;
        16'b0x1111111110x111 : cnt0=17'h4000;
        16'b111111111110x111 : cnt0=17'h8000;
        16'b0x0x0x0x0x0x1111 : cnt0=17'h400;
        16'b110x0x0x0x0x1111 : cnt0=17'h800;
        16'b10x10x0x0x0x1111 : cnt0=17'h800;
        16'b0x110x0x0x0x1111 : cnt0=17'h800;
        16'b11110x0x0x0x1111 : cnt0=17'h1000;
        16'b10x0x10x0x0x1111 : cnt0=17'h800;
        16'b0x10x10x0x0x1111 : cnt0=17'h800;
        16'b1110x10x0x0x1111 : cnt0=17'h1000;
        16'b0x0x110x0x0x1111 : cnt0=17'h800;
        16'b110x110x0x0x1111 : cnt0=17'h1000;
        16'b10x1110x0x0x1111 : cnt0=17'h1000;
        16'b0x11110x0x0x1111 : cnt0=17'h1000;
        16'b1111110x0x0x1111 : cnt0=17'h2000;
        16'b10x0x0x10x0x1111 : cnt0=17'h800;
        16'b0x10x0x10x0x1111 : cnt0=17'h800;
        16'b1110x0x10x0x1111 : cnt0=17'h1000;
        16'b0x0x10x10x0x1111 : cnt0=17'h800;
        16'b110x10x10x0x1111 : cnt0=17'h1000;
        16'b10x110x10x0x1111 : cnt0=17'h1000;
        16'b0x1110x10x0x1111 : cnt0=17'h1000;
        16'b111110x10x0x1111 : cnt0=17'h2000;
        16'b0x0x0x110x0x1111 : cnt0=17'h800;
        16'b110x0x110x0x1111 : cnt0=17'h1000;
        16'b10x10x110x0x1111 : cnt0=17'h1000;
        16'b0x110x110x0x1111 : cnt0=17'h1000;
        16'b11110x110x0x1111 : cnt0=17'h2000;
        16'b10x0x1110x0x1111 : cnt0=17'h1000;
        16'b0x10x1110x0x1111 : cnt0=17'h1000;
        16'b1110x1110x0x1111 : cnt0=17'h2000;
        16'b0x0x11110x0x1111 : cnt0=17'h1000;
        16'b110x11110x0x1111 : cnt0=17'h2000;
        16'b10x111110x0x1111 : cnt0=17'h2000;
        16'b0x1111110x0x1111 : cnt0=17'h2000;
        16'b111111110x0x1111 : cnt0=17'h4000;
        16'b10x0x0x0x10x1111 : cnt0=17'h800;
        16'b0x10x0x0x10x1111 : cnt0=17'h800;
        16'b1110x0x0x10x1111 : cnt0=17'h1000;
        16'b0x0x10x0x10x1111 : cnt0=17'h800;
        16'b110x10x0x10x1111 : cnt0=17'h1000;
        16'b10x110x0x10x1111 : cnt0=17'h1000;
        16'b0x1110x0x10x1111 : cnt0=17'h1000;
        16'b111110x0x10x1111 : cnt0=17'h2000;
        16'b0x0x0x10x10x1111 : cnt0=17'h800;
        16'b110x0x10x10x1111 : cnt0=17'h1000;
        16'b10x10x10x10x1111 : cnt0=17'h1000;
        16'b0x110x10x10x1111 : cnt0=17'h1000;
        16'b11110x10x10x1111 : cnt0=17'h2000;
        16'b10x0x110x10x1111 : cnt0=17'h1000;
        16'b0x10x110x10x1111 : cnt0=17'h1000;
        16'b1110x110x10x1111 : cnt0=17'h2000;
        16'b0x0x1110x10x1111 : cnt0=17'h1000;
        16'b110x1110x10x1111 : cnt0=17'h2000;
        16'b10x11110x10x1111 : cnt0=17'h2000;
        16'b0x111110x10x1111 : cnt0=17'h2000;
        16'b11111110x10x1111 : cnt0=17'h4000;
        16'b0x0x0x0x110x1111 : cnt0=17'h800;
        16'b110x0x0x110x1111 : cnt0=17'h1000;
        16'b10x10x0x110x1111 : cnt0=17'h1000;
        16'b0x110x0x110x1111 : cnt0=17'h1000;
        16'b11110x0x110x1111 : cnt0=17'h2000;
        16'b10x0x10x110x1111 : cnt0=17'h1000;
        16'b0x10x10x110x1111 : cnt0=17'h1000;
        16'b1110x10x110x1111 : cnt0=17'h2000;
        16'b0x0x110x110x1111 : cnt0=17'h1000;
        16'b110x110x110x1111 : cnt0=17'h2000;
        16'b10x1110x110x1111 : cnt0=17'h2000;
        16'b0x11110x110x1111 : cnt0=17'h2000;
        16'b1111110x110x1111 : cnt0=17'h4000;
        16'b10x0x0x1110x1111 : cnt0=17'h1000;
        16'b0x10x0x1110x1111 : cnt0=17'h1000;
        16'b1110x0x1110x1111 : cnt0=17'h2000;
        16'b0x0x10x1110x1111 : cnt0=17'h1000;
        16'b110x10x1110x1111 : cnt0=17'h2000;
        16'b10x110x1110x1111 : cnt0=17'h2000;
        16'b0x1110x1110x1111 : cnt0=17'h2000;
        16'b111110x1110x1111 : cnt0=17'h4000;
        16'b0x0x0x11110x1111 : cnt0=17'h1000;
        16'b110x0x11110x1111 : cnt0=17'h2000;
        16'b10x10x11110x1111 : cnt0=17'h2000;
        16'b0x110x11110x1111 : cnt0=17'h2000;
        16'b11110x11110x1111 : cnt0=17'h4000;
        16'b10x0x111110x1111 : cnt0=17'h2000;
        16'b0x10x111110x1111 : cnt0=17'h2000;
        16'b1110x111110x1111 : cnt0=17'h4000;
        16'b0x0x1111110x1111 : cnt0=17'h2000;
        16'b110x1111110x1111 : cnt0=17'h4000;
        16'b10x11111110x1111 : cnt0=17'h4000;
        16'b0x111111110x1111 : cnt0=17'h4000;
        16'b11111111110x1111 : cnt0=17'h8000;
        16'b10x0x0x0x0x11111 : cnt0=17'h800;
        16'b0x10x0x0x0x11111 : cnt0=17'h800;
        16'b1110x0x0x0x11111 : cnt0=17'h1000;
        16'b0x0x10x0x0x11111 : cnt0=17'h800;
        16'b110x10x0x0x11111 : cnt0=17'h1000;
        16'b10x110x0x0x11111 : cnt0=17'h1000;
        16'b0x1110x0x0x11111 : cnt0=17'h1000;
        16'b111110x0x0x11111 : cnt0=17'h2000;
        16'b0x0x0x10x0x11111 : cnt0=17'h800;
        16'b110x0x10x0x11111 : cnt0=17'h1000;
        16'b10x10x10x0x11111 : cnt0=17'h1000;
        16'b0x110x10x0x11111 : cnt0=17'h1000;
        16'b11110x10x0x11111 : cnt0=17'h2000;
        16'b10x0x110x0x11111 : cnt0=17'h1000;
        16'b0x10x110x0x11111 : cnt0=17'h1000;
        16'b1110x110x0x11111 : cnt0=17'h2000;
        16'b0x0x1110x0x11111 : cnt0=17'h1000;
        16'b110x1110x0x11111 : cnt0=17'h2000;
        16'b10x11110x0x11111 : cnt0=17'h2000;
        16'b0x111110x0x11111 : cnt0=17'h2000;
        16'b11111110x0x11111 : cnt0=17'h4000;
        16'b0x0x0x0x10x11111 : cnt0=17'h800;
        16'b110x0x0x10x11111 : cnt0=17'h1000;
        16'b10x10x0x10x11111 : cnt0=17'h1000;
        16'b0x110x0x10x11111 : cnt0=17'h1000;
        16'b11110x0x10x11111 : cnt0=17'h2000;
        16'b10x0x10x10x11111 : cnt0=17'h1000;
        16'b0x10x10x10x11111 : cnt0=17'h1000;
        16'b1110x10x10x11111 : cnt0=17'h2000;
        16'b0x0x110x10x11111 : cnt0=17'h1000;
        16'b110x110x10x11111 : cnt0=17'h2000;
        16'b10x1110x10x11111 : cnt0=17'h2000;
        16'b0x11110x10x11111 : cnt0=17'h2000;
        16'b1111110x10x11111 : cnt0=17'h4000;
        16'b10x0x0x110x11111 : cnt0=17'h1000;
        16'b0x10x0x110x11111 : cnt0=17'h1000;
        16'b1110x0x110x11111 : cnt0=17'h2000;
        16'b0x0x10x110x11111 : cnt0=17'h1000;
        16'b110x10x110x11111 : cnt0=17'h2000;
        16'b10x110x110x11111 : cnt0=17'h2000;
        16'b0x1110x110x11111 : cnt0=17'h2000;
        16'b111110x110x11111 : cnt0=17'h4000;
        16'b0x0x0x1110x11111 : cnt0=17'h1000;
        16'b110x0x1110x11111 : cnt0=17'h2000;
        16'b10x10x1110x11111 : cnt0=17'h2000;
        16'b0x110x1110x11111 : cnt0=17'h2000;
        16'b11110x1110x11111 : cnt0=17'h4000;
        16'b10x0x11110x11111 : cnt0=17'h2000;
        16'b0x10x11110x11111 : cnt0=17'h2000;
        16'b1110x11110x11111 : cnt0=17'h4000;
        16'b0x0x111110x11111 : cnt0=17'h2000;
        16'b110x111110x11111 : cnt0=17'h4000;
        16'b10x1111110x11111 : cnt0=17'h4000;
        16'b0x11111110x11111 : cnt0=17'h4000;
        16'b1111111110x11111 : cnt0=17'h8000;
        16'b0x0x0x0x0x111111 : cnt0=17'h800;
        16'b110x0x0x0x111111 : cnt0=17'h1000;
        16'b10x10x0x0x111111 : cnt0=17'h1000;
        16'b0x110x0x0x111111 : cnt0=17'h1000;
        16'b11110x0x0x111111 : cnt0=17'h2000;
        16'b10x0x10x0x111111 : cnt0=17'h1000;
        16'b0x10x10x0x111111 : cnt0=17'h1000;
        16'b1110x10x0x111111 : cnt0=17'h2000;
        16'b0x0x110x0x111111 : cnt0=17'h1000;
        16'b110x110x0x111111 : cnt0=17'h2000;
        16'b10x1110x0x111111 : cnt0=17'h2000;
        16'b0x11110x0x111111 : cnt0=17'h2000;
        16'b1111110x0x111111 : cnt0=17'h4000;
        16'b10x0x0x10x111111 : cnt0=17'h1000;
        16'b0x10x0x10x111111 : cnt0=17'h1000;
        16'b1110x0x10x111111 : cnt0=17'h2000;
        16'b0x0x10x10x111111 : cnt0=17'h1000;
        16'b110x10x10x111111 : cnt0=17'h2000;
        16'b10x110x10x111111 : cnt0=17'h2000;
        16'b0x1110x10x111111 : cnt0=17'h2000;
        16'b111110x10x111111 : cnt0=17'h4000;
        16'b0x0x0x110x111111 : cnt0=17'h1000;
        16'b110x0x110x111111 : cnt0=17'h2000;
        16'b10x10x110x111111 : cnt0=17'h2000;
        16'b0x110x110x111111 : cnt0=17'h2000;
        16'b11110x110x111111 : cnt0=17'h4000;
        16'b10x0x1110x111111 : cnt0=17'h2000;
        16'b0x10x1110x111111 : cnt0=17'h2000;
        16'b1110x1110x111111 : cnt0=17'h4000;
        16'b0x0x11110x111111 : cnt0=17'h2000;
        16'b110x11110x111111 : cnt0=17'h4000;
        16'b10x111110x111111 : cnt0=17'h4000;
        16'b0x1111110x111111 : cnt0=17'h4000;
        16'b111111110x111111 : cnt0=17'h8000;
        16'b10x0x0x0x1111111 : cnt0=17'h1000;
        16'b0x10x0x0x1111111 : cnt0=17'h1000;
        16'b1110x0x0x1111111 : cnt0=17'h2000;
        16'b0x0x10x0x1111111 : cnt0=17'h1000;
        16'b110x10x0x1111111 : cnt0=17'h2000;
        16'b10x110x0x1111111 : cnt0=17'h2000;
        16'b0x1110x0x1111111 : cnt0=17'h2000;
        16'b111110x0x1111111 : cnt0=17'h4000;
        16'b0x0x0x10x1111111 : cnt0=17'h1000;
        16'b110x0x10x1111111 : cnt0=17'h2000;
        16'b10x10x10x1111111 : cnt0=17'h2000;
        16'b0x110x10x1111111 : cnt0=17'h2000;
        16'b11110x10x1111111 : cnt0=17'h4000;
        16'b10x0x110x1111111 : cnt0=17'h2000;
        16'b0x10x110x1111111 : cnt0=17'h2000;
        16'b1110x110x1111111 : cnt0=17'h4000;
        16'b0x0x1110x1111111 : cnt0=17'h2000;
        16'b110x1110x1111111 : cnt0=17'h4000;
        16'b10x11110x1111111 : cnt0=17'h4000;
        16'b0x111110x1111111 : cnt0=17'h4000;
        16'b11111110x1111111 : cnt0=17'h8000;
        16'b0x0x0x0x11111111 : cnt0=17'h1000;
        16'b110x0x0x11111111 : cnt0=17'h2000;
        16'b10x10x0x11111111 : cnt0=17'h2000;
        16'b0x110x0x11111111 : cnt0=17'h2000;
        16'b11110x0x11111111 : cnt0=17'h4000;
        16'b10x0x10x11111111 : cnt0=17'h2000;
        16'b0x10x10x11111111 : cnt0=17'h2000;
        16'b1110x10x11111111 : cnt0=17'h4000;
        16'b0x0x110x11111111 : cnt0=17'h2000;
        16'b110x110x11111111 : cnt0=17'h4000;
        16'b10x1110x11111111 : cnt0=17'h4000;
        16'b0x11110x11111111 : cnt0=17'h4000;
        16'b1111110x11111111 : cnt0=17'h8000;
        16'b10x0x0x111111111 : cnt0=17'h2000;
        16'b0x10x0x111111111 : cnt0=17'h2000;
        16'b1110x0x111111111 : cnt0=17'h4000;
        16'b0x0x10x111111111 : cnt0=17'h2000;
        16'b110x10x111111111 : cnt0=17'h4000;
        16'b10x110x111111111 : cnt0=17'h4000;
        16'b0x1110x111111111 : cnt0=17'h4000;
        16'b111110x111111111 : cnt0=17'h8000;
        16'b0x0x0x1111111111 : cnt0=17'h2000;
        16'b110x0x1111111111 : cnt0=17'h4000;
        16'b10x10x1111111111 : cnt0=17'h4000;
        16'b0x110x1111111111 : cnt0=17'h4000;
        16'b11110x1111111111 : cnt0=17'h8000;
        16'b10x0x11111111111 : cnt0=17'h4000;
        16'b0x10x11111111111 : cnt0=17'h4000;
        16'b1110x11111111111 : cnt0=17'h8000;
        16'b0x0x111111111111 : cnt0=17'h4000;
        16'b110x111111111111 : cnt0=17'h8000;
        16'b10x1111111111111 : cnt0=17'h8000;
        16'b0x11111111111111 : cnt0=17'h8000;
        16'b1111111111111111 : cnt0=17'h10000;
    endcase

  endfunction
  function [0:0] tail0;
    input [15:0] bits;
    casex(bits)
        16'b0x0x0x0x0x0x0x0x : tail0=1'b0;
        16'b10x0x0x0x0x0x0x0 : tail0=1'b0;
        16'b110x0x0x0x0x0x0x : tail0=1'b0;
        16'b0x10x0x0x0x0x0x0 : tail0=1'b0;
        16'b1110x0x0x0x0x0x0 : tail0=1'b0;
        16'b10x10x0x0x0x0x0x : tail0=1'b0;
        16'b0x110x0x0x0x0x0x : tail0=1'b0;
        16'b11110x0x0x0x0x0x : tail0=1'b0;
        16'b0x0x10x0x0x0x0x0 : tail0=1'b0;
        16'b110x10x0x0x0x0x0 : tail0=1'b0;
        16'b10x110x0x0x0x0x0 : tail0=1'b0;
        16'b0x1110x0x0x0x0x0 : tail0=1'b0;
        16'b111110x0x0x0x0x0 : tail0=1'b0;
        16'b10x0x10x0x0x0x0x : tail0=1'b0;
        16'b0x10x10x0x0x0x0x : tail0=1'b0;
        16'b1110x10x0x0x0x0x : tail0=1'b0;
        16'b0x0x110x0x0x0x0x : tail0=1'b0;
        16'b110x110x0x0x0x0x : tail0=1'b0;
        16'b10x1110x0x0x0x0x : tail0=1'b0;
        16'b0x11110x0x0x0x0x : tail0=1'b0;
        16'b1111110x0x0x0x0x : tail0=1'b0;
        16'b0x0x0x10x0x0x0x0 : tail0=1'b0;
        16'b110x0x10x0x0x0x0 : tail0=1'b0;
        16'b10x10x10x0x0x0x0 : tail0=1'b0;
        16'b0x110x10x0x0x0x0 : tail0=1'b0;
        16'b11110x10x0x0x0x0 : tail0=1'b0;
        16'b10x0x110x0x0x0x0 : tail0=1'b0;
        16'b0x10x110x0x0x0x0 : tail0=1'b0;
        16'b1110x110x0x0x0x0 : tail0=1'b0;
        16'b0x0x1110x0x0x0x0 : tail0=1'b0;
        16'b110x1110x0x0x0x0 : tail0=1'b0;
        16'b10x11110x0x0x0x0 : tail0=1'b0;
        16'b0x111110x0x0x0x0 : tail0=1'b0;
        16'b11111110x0x0x0x0 : tail0=1'b0;
        16'b10x0x0x10x0x0x0x : tail0=1'b0;
        16'b0x10x0x10x0x0x0x : tail0=1'b0;
        16'b1110x0x10x0x0x0x : tail0=1'b0;
        16'b0x0x10x10x0x0x0x : tail0=1'b0;
        16'b110x10x10x0x0x0x : tail0=1'b0;
        16'b10x110x10x0x0x0x : tail0=1'b0;
        16'b0x1110x10x0x0x0x : tail0=1'b0;
        16'b111110x10x0x0x0x : tail0=1'b0;
        16'b0x0x0x110x0x0x0x : tail0=1'b0;
        16'b110x0x110x0x0x0x : tail0=1'b0;
        16'b10x10x110x0x0x0x : tail0=1'b0;
        16'b0x110x110x0x0x0x : tail0=1'b0;
        16'b11110x110x0x0x0x : tail0=1'b0;
        16'b10x0x1110x0x0x0x : tail0=1'b0;
        16'b0x10x1110x0x0x0x : tail0=1'b0;
        16'b1110x1110x0x0x0x : tail0=1'b0;
        16'b0x0x11110x0x0x0x : tail0=1'b0;
        16'b110x11110x0x0x0x : tail0=1'b0;
        16'b10x111110x0x0x0x : tail0=1'b0;
        16'b0x1111110x0x0x0x : tail0=1'b0;
        16'b111111110x0x0x0x : tail0=1'b0;
        16'b0x0x0x0x10x0x0x0 : tail0=1'b0;
        16'b110x0x0x10x0x0x0 : tail0=1'b0;
        16'b10x10x0x10x0x0x0 : tail0=1'b0;
        16'b0x110x0x10x0x0x0 : tail0=1'b0;
        16'b11110x0x10x0x0x0 : tail0=1'b0;
        16'b10x0x10x10x0x0x0 : tail0=1'b0;
        16'b0x10x10x10x0x0x0 : tail0=1'b0;
        16'b1110x10x10x0x0x0 : tail0=1'b0;
        16'b0x0x110x10x0x0x0 : tail0=1'b0;
        16'b110x110x10x0x0x0 : tail0=1'b0;
        16'b10x1110x10x0x0x0 : tail0=1'b0;
        16'b0x11110x10x0x0x0 : tail0=1'b0;
        16'b1111110x10x0x0x0 : tail0=1'b0;
        16'b10x0x0x110x0x0x0 : tail0=1'b0;
        16'b0x10x0x110x0x0x0 : tail0=1'b0;
        16'b1110x0x110x0x0x0 : tail0=1'b0;
        16'b0x0x10x110x0x0x0 : tail0=1'b0;
        16'b110x10x110x0x0x0 : tail0=1'b0;
        16'b10x110x110x0x0x0 : tail0=1'b0;
        16'b0x1110x110x0x0x0 : tail0=1'b0;
        16'b111110x110x0x0x0 : tail0=1'b0;
        16'b0x0x0x1110x0x0x0 : tail0=1'b0;
        16'b110x0x1110x0x0x0 : tail0=1'b0;
        16'b10x10x1110x0x0x0 : tail0=1'b0;
        16'b0x110x1110x0x0x0 : tail0=1'b0;
        16'b11110x1110x0x0x0 : tail0=1'b0;
        16'b10x0x11110x0x0x0 : tail0=1'b0;
        16'b0x10x11110x0x0x0 : tail0=1'b0;
        16'b1110x11110x0x0x0 : tail0=1'b0;
        16'b0x0x111110x0x0x0 : tail0=1'b0;
        16'b110x111110x0x0x0 : tail0=1'b0;
        16'b10x1111110x0x0x0 : tail0=1'b0;
        16'b0x11111110x0x0x0 : tail0=1'b0;
        16'b1111111110x0x0x0 : tail0=1'b0;
        16'b10x0x0x0x10x0x0x : tail0=1'b0;
        16'b0x10x0x0x10x0x0x : tail0=1'b0;
        16'b1110x0x0x10x0x0x : tail0=1'b0;
        16'b0x0x10x0x10x0x0x : tail0=1'b0;
        16'b110x10x0x10x0x0x : tail0=1'b0;
        16'b10x110x0x10x0x0x : tail0=1'b0;
        16'b0x1110x0x10x0x0x : tail0=1'b0;
        16'b111110x0x10x0x0x : tail0=1'b0;
        16'b0x0x0x10x10x0x0x : tail0=1'b0;
        16'b110x0x10x10x0x0x : tail0=1'b0;
        16'b10x10x10x10x0x0x : tail0=1'b0;
        16'b0x110x10x10x0x0x : tail0=1'b0;
        16'b11110x10x10x0x0x : tail0=1'b0;
        16'b10x0x110x10x0x0x : tail0=1'b0;
        16'b0x10x110x10x0x0x : tail0=1'b0;
        16'b1110x110x10x0x0x : tail0=1'b0;
        16'b0x0x1110x10x0x0x : tail0=1'b0;
        16'b110x1110x10x0x0x : tail0=1'b0;
        16'b10x11110x10x0x0x : tail0=1'b0;
        16'b0x111110x10x0x0x : tail0=1'b0;
        16'b11111110x10x0x0x : tail0=1'b0;
        16'b0x0x0x0x110x0x0x : tail0=1'b0;
        16'b110x0x0x110x0x0x : tail0=1'b0;
        16'b10x10x0x110x0x0x : tail0=1'b0;
        16'b0x110x0x110x0x0x : tail0=1'b0;
        16'b11110x0x110x0x0x : tail0=1'b0;
        16'b10x0x10x110x0x0x : tail0=1'b0;
        16'b0x10x10x110x0x0x : tail0=1'b0;
        16'b1110x10x110x0x0x : tail0=1'b0;
        16'b0x0x110x110x0x0x : tail0=1'b0;
        16'b110x110x110x0x0x : tail0=1'b0;
        16'b10x1110x110x0x0x : tail0=1'b0;
        16'b0x11110x110x0x0x : tail0=1'b0;
        16'b1111110x110x0x0x : tail0=1'b0;
        16'b10x0x0x1110x0x0x : tail0=1'b0;
        16'b0x10x0x1110x0x0x : tail0=1'b0;
        16'b1110x0x1110x0x0x : tail0=1'b0;
        16'b0x0x10x1110x0x0x : tail0=1'b0;
        16'b110x10x1110x0x0x : tail0=1'b0;
        16'b10x110x1110x0x0x : tail0=1'b0;
        16'b0x1110x1110x0x0x : tail0=1'b0;
        16'b111110x1110x0x0x : tail0=1'b0;
        16'b0x0x0x11110x0x0x : tail0=1'b0;
        16'b110x0x11110x0x0x : tail0=1'b0;
        16'b10x10x11110x0x0x : tail0=1'b0;
        16'b0x110x11110x0x0x : tail0=1'b0;
        16'b11110x11110x0x0x : tail0=1'b0;
        16'b10x0x111110x0x0x : tail0=1'b0;
        16'b0x10x111110x0x0x : tail0=1'b0;
        16'b1110x111110x0x0x : tail0=1'b0;
        16'b0x0x1111110x0x0x : tail0=1'b0;
        16'b110x1111110x0x0x : tail0=1'b0;
        16'b10x11111110x0x0x : tail0=1'b0;
        16'b0x111111110x0x0x : tail0=1'b0;
        16'b11111111110x0x0x : tail0=1'b0;
        16'b0x0x0x0x0x10x0x0 : tail0=1'b0;
        16'b110x0x0x0x10x0x0 : tail0=1'b0;
        16'b10x10x0x0x10x0x0 : tail0=1'b0;
        16'b0x110x0x0x10x0x0 : tail0=1'b0;
        16'b11110x0x0x10x0x0 : tail0=1'b0;
        16'b10x0x10x0x10x0x0 : tail0=1'b0;
        16'b0x10x10x0x10x0x0 : tail0=1'b0;
        16'b1110x10x0x10x0x0 : tail0=1'b0;
        16'b0x0x110x0x10x0x0 : tail0=1'b0;
        16'b110x110x0x10x0x0 : tail0=1'b0;
        16'b10x1110x0x10x0x0 : tail0=1'b0;
        16'b0x11110x0x10x0x0 : tail0=1'b0;
        16'b1111110x0x10x0x0 : tail0=1'b0;
        16'b10x0x0x10x10x0x0 : tail0=1'b0;
        16'b0x10x0x10x10x0x0 : tail0=1'b0;
        16'b1110x0x10x10x0x0 : tail0=1'b0;
        16'b0x0x10x10x10x0x0 : tail0=1'b0;
        16'b110x10x10x10x0x0 : tail0=1'b0;
        16'b10x110x10x10x0x0 : tail0=1'b0;
        16'b0x1110x10x10x0x0 : tail0=1'b0;
        16'b111110x10x10x0x0 : tail0=1'b0;
        16'b0x0x0x110x10x0x0 : tail0=1'b0;
        16'b110x0x110x10x0x0 : tail0=1'b0;
        16'b10x10x110x10x0x0 : tail0=1'b0;
        16'b0x110x110x10x0x0 : tail0=1'b0;
        16'b11110x110x10x0x0 : tail0=1'b0;
        16'b10x0x1110x10x0x0 : tail0=1'b0;
        16'b0x10x1110x10x0x0 : tail0=1'b0;
        16'b1110x1110x10x0x0 : tail0=1'b0;
        16'b0x0x11110x10x0x0 : tail0=1'b0;
        16'b110x11110x10x0x0 : tail0=1'b0;
        16'b10x111110x10x0x0 : tail0=1'b0;
        16'b0x1111110x10x0x0 : tail0=1'b0;
        16'b111111110x10x0x0 : tail0=1'b0;
        16'b10x0x0x0x110x0x0 : tail0=1'b0;
        16'b0x10x0x0x110x0x0 : tail0=1'b0;
        16'b1110x0x0x110x0x0 : tail0=1'b0;
        16'b0x0x10x0x110x0x0 : tail0=1'b0;
        16'b110x10x0x110x0x0 : tail0=1'b0;
        16'b10x110x0x110x0x0 : tail0=1'b0;
        16'b0x1110x0x110x0x0 : tail0=1'b0;
        16'b111110x0x110x0x0 : tail0=1'b0;
        16'b0x0x0x10x110x0x0 : tail0=1'b0;
        16'b110x0x10x110x0x0 : tail0=1'b0;
        16'b10x10x10x110x0x0 : tail0=1'b0;
        16'b0x110x10x110x0x0 : tail0=1'b0;
        16'b11110x10x110x0x0 : tail0=1'b0;
        16'b10x0x110x110x0x0 : tail0=1'b0;
        16'b0x10x110x110x0x0 : tail0=1'b0;
        16'b1110x110x110x0x0 : tail0=1'b0;
        16'b0x0x1110x110x0x0 : tail0=1'b0;
        16'b110x1110x110x0x0 : tail0=1'b0;
        16'b10x11110x110x0x0 : tail0=1'b0;
        16'b0x111110x110x0x0 : tail0=1'b0;
        16'b11111110x110x0x0 : tail0=1'b0;
        16'b0x0x0x0x1110x0x0 : tail0=1'b0;
        16'b110x0x0x1110x0x0 : tail0=1'b0;
        16'b10x10x0x1110x0x0 : tail0=1'b0;
        16'b0x110x0x1110x0x0 : tail0=1'b0;
        16'b11110x0x1110x0x0 : tail0=1'b0;
        16'b10x0x10x1110x0x0 : tail0=1'b0;
        16'b0x10x10x1110x0x0 : tail0=1'b0;
        16'b1110x10x1110x0x0 : tail0=1'b0;
        16'b0x0x110x1110x0x0 : tail0=1'b0;
        16'b110x110x1110x0x0 : tail0=1'b0;
        16'b10x1110x1110x0x0 : tail0=1'b0;
        16'b0x11110x1110x0x0 : tail0=1'b0;
        16'b1111110x1110x0x0 : tail0=1'b0;
        16'b10x0x0x11110x0x0 : tail0=1'b0;
        16'b0x10x0x11110x0x0 : tail0=1'b0;
        16'b1110x0x11110x0x0 : tail0=1'b0;
        16'b0x0x10x11110x0x0 : tail0=1'b0;
        16'b110x10x11110x0x0 : tail0=1'b0;
        16'b10x110x11110x0x0 : tail0=1'b0;
        16'b0x1110x11110x0x0 : tail0=1'b0;
        16'b111110x11110x0x0 : tail0=1'b0;
        16'b0x0x0x111110x0x0 : tail0=1'b0;
        16'b110x0x111110x0x0 : tail0=1'b0;
        16'b10x10x111110x0x0 : tail0=1'b0;
        16'b0x110x111110x0x0 : tail0=1'b0;
        16'b11110x111110x0x0 : tail0=1'b0;
        16'b10x0x1111110x0x0 : tail0=1'b0;
        16'b0x10x1111110x0x0 : tail0=1'b0;
        16'b1110x1111110x0x0 : tail0=1'b0;
        16'b0x0x11111110x0x0 : tail0=1'b0;
        16'b110x11111110x0x0 : tail0=1'b0;
        16'b10x111111110x0x0 : tail0=1'b0;
        16'b0x1111111110x0x0 : tail0=1'b0;
        16'b111111111110x0x0 : tail0=1'b0;
        16'b10x0x0x0x0x10x0x : tail0=1'b0;
        16'b0x10x0x0x0x10x0x : tail0=1'b0;
        16'b1110x0x0x0x10x0x : tail0=1'b0;
        16'b0x0x10x0x0x10x0x : tail0=1'b0;
        16'b110x10x0x0x10x0x : tail0=1'b0;
        16'b10x110x0x0x10x0x : tail0=1'b0;
        16'b0x1110x0x0x10x0x : tail0=1'b0;
        16'b111110x0x0x10x0x : tail0=1'b0;
        16'b0x0x0x10x0x10x0x : tail0=1'b0;
        16'b110x0x10x0x10x0x : tail0=1'b0;
        16'b10x10x10x0x10x0x : tail0=1'b0;
        16'b0x110x10x0x10x0x : tail0=1'b0;
        16'b11110x10x0x10x0x : tail0=1'b0;
        16'b10x0x110x0x10x0x : tail0=1'b0;
        16'b0x10x110x0x10x0x : tail0=1'b0;
        16'b1110x110x0x10x0x : tail0=1'b0;
        16'b0x0x1110x0x10x0x : tail0=1'b0;
        16'b110x1110x0x10x0x : tail0=1'b0;
        16'b10x11110x0x10x0x : tail0=1'b0;
        16'b0x111110x0x10x0x : tail0=1'b0;
        16'b11111110x0x10x0x : tail0=1'b0;
        16'b0x0x0x0x10x10x0x : tail0=1'b0;
        16'b110x0x0x10x10x0x : tail0=1'b0;
        16'b10x10x0x10x10x0x : tail0=1'b0;
        16'b0x110x0x10x10x0x : tail0=1'b0;
        16'b11110x0x10x10x0x : tail0=1'b0;
        16'b10x0x10x10x10x0x : tail0=1'b0;
        16'b0x10x10x10x10x0x : tail0=1'b0;
        16'b1110x10x10x10x0x : tail0=1'b0;
        16'b0x0x110x10x10x0x : tail0=1'b0;
        16'b110x110x10x10x0x : tail0=1'b0;
        16'b10x1110x10x10x0x : tail0=1'b0;
        16'b0x11110x10x10x0x : tail0=1'b0;
        16'b1111110x10x10x0x : tail0=1'b0;
        16'b10x0x0x110x10x0x : tail0=1'b0;
        16'b0x10x0x110x10x0x : tail0=1'b0;
        16'b1110x0x110x10x0x : tail0=1'b0;
        16'b0x0x10x110x10x0x : tail0=1'b0;
        16'b110x10x110x10x0x : tail0=1'b0;
        16'b10x110x110x10x0x : tail0=1'b0;
        16'b0x1110x110x10x0x : tail0=1'b0;
        16'b111110x110x10x0x : tail0=1'b0;
        16'b0x0x0x1110x10x0x : tail0=1'b0;
        16'b110x0x1110x10x0x : tail0=1'b0;
        16'b10x10x1110x10x0x : tail0=1'b0;
        16'b0x110x1110x10x0x : tail0=1'b0;
        16'b11110x1110x10x0x : tail0=1'b0;
        16'b10x0x11110x10x0x : tail0=1'b0;
        16'b0x10x11110x10x0x : tail0=1'b0;
        16'b1110x11110x10x0x : tail0=1'b0;
        16'b0x0x111110x10x0x : tail0=1'b0;
        16'b110x111110x10x0x : tail0=1'b0;
        16'b10x1111110x10x0x : tail0=1'b0;
        16'b0x11111110x10x0x : tail0=1'b0;
        16'b1111111110x10x0x : tail0=1'b0;
        16'b0x0x0x0x0x110x0x : tail0=1'b0;
        16'b110x0x0x0x110x0x : tail0=1'b0;
        16'b10x10x0x0x110x0x : tail0=1'b0;
        16'b0x110x0x0x110x0x : tail0=1'b0;
        16'b11110x0x0x110x0x : tail0=1'b0;
        16'b10x0x10x0x110x0x : tail0=1'b0;
        16'b0x10x10x0x110x0x : tail0=1'b0;
        16'b1110x10x0x110x0x : tail0=1'b0;
        16'b0x0x110x0x110x0x : tail0=1'b0;
        16'b110x110x0x110x0x : tail0=1'b0;
        16'b10x1110x0x110x0x : tail0=1'b0;
        16'b0x11110x0x110x0x : tail0=1'b0;
        16'b1111110x0x110x0x : tail0=1'b0;
        16'b10x0x0x10x110x0x : tail0=1'b0;
        16'b0x10x0x10x110x0x : tail0=1'b0;
        16'b1110x0x10x110x0x : tail0=1'b0;
        16'b0x0x10x10x110x0x : tail0=1'b0;
        16'b110x10x10x110x0x : tail0=1'b0;
        16'b10x110x10x110x0x : tail0=1'b0;
        16'b0x1110x10x110x0x : tail0=1'b0;
        16'b111110x10x110x0x : tail0=1'b0;
        16'b0x0x0x110x110x0x : tail0=1'b0;
        16'b110x0x110x110x0x : tail0=1'b0;
        16'b10x10x110x110x0x : tail0=1'b0;
        16'b0x110x110x110x0x : tail0=1'b0;
        16'b11110x110x110x0x : tail0=1'b0;
        16'b10x0x1110x110x0x : tail0=1'b0;
        16'b0x10x1110x110x0x : tail0=1'b0;
        16'b1110x1110x110x0x : tail0=1'b0;
        16'b0x0x11110x110x0x : tail0=1'b0;
        16'b110x11110x110x0x : tail0=1'b0;
        16'b10x111110x110x0x : tail0=1'b0;
        16'b0x1111110x110x0x : tail0=1'b0;
        16'b111111110x110x0x : tail0=1'b0;
        16'b10x0x0x0x1110x0x : tail0=1'b0;
        16'b0x10x0x0x1110x0x : tail0=1'b0;
        16'b1110x0x0x1110x0x : tail0=1'b0;
        16'b0x0x10x0x1110x0x : tail0=1'b0;
        16'b110x10x0x1110x0x : tail0=1'b0;
        16'b10x110x0x1110x0x : tail0=1'b0;
        16'b0x1110x0x1110x0x : tail0=1'b0;
        16'b111110x0x1110x0x : tail0=1'b0;
        16'b0x0x0x10x1110x0x : tail0=1'b0;
        16'b110x0x10x1110x0x : tail0=1'b0;
        16'b10x10x10x1110x0x : tail0=1'b0;
        16'b0x110x10x1110x0x : tail0=1'b0;
        16'b11110x10x1110x0x : tail0=1'b0;
        16'b10x0x110x1110x0x : tail0=1'b0;
        16'b0x10x110x1110x0x : tail0=1'b0;
        16'b1110x110x1110x0x : tail0=1'b0;
        16'b0x0x1110x1110x0x : tail0=1'b0;
        16'b110x1110x1110x0x : tail0=1'b0;
        16'b10x11110x1110x0x : tail0=1'b0;
        16'b0x111110x1110x0x : tail0=1'b0;
        16'b11111110x1110x0x : tail0=1'b0;
        16'b0x0x0x0x11110x0x : tail0=1'b0;
        16'b110x0x0x11110x0x : tail0=1'b0;
        16'b10x10x0x11110x0x : tail0=1'b0;
        16'b0x110x0x11110x0x : tail0=1'b0;
        16'b11110x0x11110x0x : tail0=1'b0;
        16'b10x0x10x11110x0x : tail0=1'b0;
        16'b0x10x10x11110x0x : tail0=1'b0;
        16'b1110x10x11110x0x : tail0=1'b0;
        16'b0x0x110x11110x0x : tail0=1'b0;
        16'b110x110x11110x0x : tail0=1'b0;
        16'b10x1110x11110x0x : tail0=1'b0;
        16'b0x11110x11110x0x : tail0=1'b0;
        16'b1111110x11110x0x : tail0=1'b0;
        16'b10x0x0x111110x0x : tail0=1'b0;
        16'b0x10x0x111110x0x : tail0=1'b0;
        16'b1110x0x111110x0x : tail0=1'b0;
        16'b0x0x10x111110x0x : tail0=1'b0;
        16'b110x10x111110x0x : tail0=1'b0;
        16'b10x110x111110x0x : tail0=1'b0;
        16'b0x1110x111110x0x : tail0=1'b0;
        16'b111110x111110x0x : tail0=1'b0;
        16'b0x0x0x1111110x0x : tail0=1'b0;
        16'b110x0x1111110x0x : tail0=1'b0;
        16'b10x10x1111110x0x : tail0=1'b0;
        16'b0x110x1111110x0x : tail0=1'b0;
        16'b11110x1111110x0x : tail0=1'b0;
        16'b10x0x11111110x0x : tail0=1'b0;
        16'b0x10x11111110x0x : tail0=1'b0;
        16'b1110x11111110x0x : tail0=1'b0;
        16'b0x0x111111110x0x : tail0=1'b0;
        16'b110x111111110x0x : tail0=1'b0;
        16'b10x1111111110x0x : tail0=1'b0;
        16'b0x11111111110x0x : tail0=1'b0;
        16'b1111111111110x0x : tail0=1'b0;
        16'b0x0x0x0x0x0x10x0 : tail0=1'b0;
        16'b110x0x0x0x0x10x0 : tail0=1'b0;
        16'b10x10x0x0x0x10x0 : tail0=1'b0;
        16'b0x110x0x0x0x10x0 : tail0=1'b0;
        16'b11110x0x0x0x10x0 : tail0=1'b0;
        16'b10x0x10x0x0x10x0 : tail0=1'b0;
        16'b0x10x10x0x0x10x0 : tail0=1'b0;
        16'b1110x10x0x0x10x0 : tail0=1'b0;
        16'b0x0x110x0x0x10x0 : tail0=1'b0;
        16'b110x110x0x0x10x0 : tail0=1'b0;
        16'b10x1110x0x0x10x0 : tail0=1'b0;
        16'b0x11110x0x0x10x0 : tail0=1'b0;
        16'b1111110x0x0x10x0 : tail0=1'b0;
        16'b10x0x0x10x0x10x0 : tail0=1'b0;
        16'b0x10x0x10x0x10x0 : tail0=1'b0;
        16'b1110x0x10x0x10x0 : tail0=1'b0;
        16'b0x0x10x10x0x10x0 : tail0=1'b0;
        16'b110x10x10x0x10x0 : tail0=1'b0;
        16'b10x110x10x0x10x0 : tail0=1'b0;
        16'b0x1110x10x0x10x0 : tail0=1'b0;
        16'b111110x10x0x10x0 : tail0=1'b0;
        16'b0x0x0x110x0x10x0 : tail0=1'b0;
        16'b110x0x110x0x10x0 : tail0=1'b0;
        16'b10x10x110x0x10x0 : tail0=1'b0;
        16'b0x110x110x0x10x0 : tail0=1'b0;
        16'b11110x110x0x10x0 : tail0=1'b0;
        16'b10x0x1110x0x10x0 : tail0=1'b0;
        16'b0x10x1110x0x10x0 : tail0=1'b0;
        16'b1110x1110x0x10x0 : tail0=1'b0;
        16'b0x0x11110x0x10x0 : tail0=1'b0;
        16'b110x11110x0x10x0 : tail0=1'b0;
        16'b10x111110x0x10x0 : tail0=1'b0;
        16'b0x1111110x0x10x0 : tail0=1'b0;
        16'b111111110x0x10x0 : tail0=1'b0;
        16'b10x0x0x0x10x10x0 : tail0=1'b0;
        16'b0x10x0x0x10x10x0 : tail0=1'b0;
        16'b1110x0x0x10x10x0 : tail0=1'b0;
        16'b0x0x10x0x10x10x0 : tail0=1'b0;
        16'b110x10x0x10x10x0 : tail0=1'b0;
        16'b10x110x0x10x10x0 : tail0=1'b0;
        16'b0x1110x0x10x10x0 : tail0=1'b0;
        16'b111110x0x10x10x0 : tail0=1'b0;
        16'b0x0x0x10x10x10x0 : tail0=1'b0;
        16'b110x0x10x10x10x0 : tail0=1'b0;
        16'b10x10x10x10x10x0 : tail0=1'b0;
        16'b0x110x10x10x10x0 : tail0=1'b0;
        16'b11110x10x10x10x0 : tail0=1'b0;
        16'b10x0x110x10x10x0 : tail0=1'b0;
        16'b0x10x110x10x10x0 : tail0=1'b0;
        16'b1110x110x10x10x0 : tail0=1'b0;
        16'b0x0x1110x10x10x0 : tail0=1'b0;
        16'b110x1110x10x10x0 : tail0=1'b0;
        16'b10x11110x10x10x0 : tail0=1'b0;
        16'b0x111110x10x10x0 : tail0=1'b0;
        16'b11111110x10x10x0 : tail0=1'b0;
        16'b0x0x0x0x110x10x0 : tail0=1'b0;
        16'b110x0x0x110x10x0 : tail0=1'b0;
        16'b10x10x0x110x10x0 : tail0=1'b0;
        16'b0x110x0x110x10x0 : tail0=1'b0;
        16'b11110x0x110x10x0 : tail0=1'b0;
        16'b10x0x10x110x10x0 : tail0=1'b0;
        16'b0x10x10x110x10x0 : tail0=1'b0;
        16'b1110x10x110x10x0 : tail0=1'b0;
        16'b0x0x110x110x10x0 : tail0=1'b0;
        16'b110x110x110x10x0 : tail0=1'b0;
        16'b10x1110x110x10x0 : tail0=1'b0;
        16'b0x11110x110x10x0 : tail0=1'b0;
        16'b1111110x110x10x0 : tail0=1'b0;
        16'b10x0x0x1110x10x0 : tail0=1'b0;
        16'b0x10x0x1110x10x0 : tail0=1'b0;
        16'b1110x0x1110x10x0 : tail0=1'b0;
        16'b0x0x10x1110x10x0 : tail0=1'b0;
        16'b110x10x1110x10x0 : tail0=1'b0;
        16'b10x110x1110x10x0 : tail0=1'b0;
        16'b0x1110x1110x10x0 : tail0=1'b0;
        16'b111110x1110x10x0 : tail0=1'b0;
        16'b0x0x0x11110x10x0 : tail0=1'b0;
        16'b110x0x11110x10x0 : tail0=1'b0;
        16'b10x10x11110x10x0 : tail0=1'b0;
        16'b0x110x11110x10x0 : tail0=1'b0;
        16'b11110x11110x10x0 : tail0=1'b0;
        16'b10x0x111110x10x0 : tail0=1'b0;
        16'b0x10x111110x10x0 : tail0=1'b0;
        16'b1110x111110x10x0 : tail0=1'b0;
        16'b0x0x1111110x10x0 : tail0=1'b0;
        16'b110x1111110x10x0 : tail0=1'b0;
        16'b10x11111110x10x0 : tail0=1'b0;
        16'b0x111111110x10x0 : tail0=1'b0;
        16'b11111111110x10x0 : tail0=1'b0;
        16'b10x0x0x0x0x110x0 : tail0=1'b0;
        16'b0x10x0x0x0x110x0 : tail0=1'b0;
        16'b1110x0x0x0x110x0 : tail0=1'b0;
        16'b0x0x10x0x0x110x0 : tail0=1'b0;
        16'b110x10x0x0x110x0 : tail0=1'b0;
        16'b10x110x0x0x110x0 : tail0=1'b0;
        16'b0x1110x0x0x110x0 : tail0=1'b0;
        16'b111110x0x0x110x0 : tail0=1'b0;
        16'b0x0x0x10x0x110x0 : tail0=1'b0;
        16'b110x0x10x0x110x0 : tail0=1'b0;
        16'b10x10x10x0x110x0 : tail0=1'b0;
        16'b0x110x10x0x110x0 : tail0=1'b0;
        16'b11110x10x0x110x0 : tail0=1'b0;
        16'b10x0x110x0x110x0 : tail0=1'b0;
        16'b0x10x110x0x110x0 : tail0=1'b0;
        16'b1110x110x0x110x0 : tail0=1'b0;
        16'b0x0x1110x0x110x0 : tail0=1'b0;
        16'b110x1110x0x110x0 : tail0=1'b0;
        16'b10x11110x0x110x0 : tail0=1'b0;
        16'b0x111110x0x110x0 : tail0=1'b0;
        16'b11111110x0x110x0 : tail0=1'b0;
        16'b0x0x0x0x10x110x0 : tail0=1'b0;
        16'b110x0x0x10x110x0 : tail0=1'b0;
        16'b10x10x0x10x110x0 : tail0=1'b0;
        16'b0x110x0x10x110x0 : tail0=1'b0;
        16'b11110x0x10x110x0 : tail0=1'b0;
        16'b10x0x10x10x110x0 : tail0=1'b0;
        16'b0x10x10x10x110x0 : tail0=1'b0;
        16'b1110x10x10x110x0 : tail0=1'b0;
        16'b0x0x110x10x110x0 : tail0=1'b0;
        16'b110x110x10x110x0 : tail0=1'b0;
        16'b10x1110x10x110x0 : tail0=1'b0;
        16'b0x11110x10x110x0 : tail0=1'b0;
        16'b1111110x10x110x0 : tail0=1'b0;
        16'b10x0x0x110x110x0 : tail0=1'b0;
        16'b0x10x0x110x110x0 : tail0=1'b0;
        16'b1110x0x110x110x0 : tail0=1'b0;
        16'b0x0x10x110x110x0 : tail0=1'b0;
        16'b110x10x110x110x0 : tail0=1'b0;
        16'b10x110x110x110x0 : tail0=1'b0;
        16'b0x1110x110x110x0 : tail0=1'b0;
        16'b111110x110x110x0 : tail0=1'b0;
        16'b0x0x0x1110x110x0 : tail0=1'b0;
        16'b110x0x1110x110x0 : tail0=1'b0;
        16'b10x10x1110x110x0 : tail0=1'b0;
        16'b0x110x1110x110x0 : tail0=1'b0;
        16'b11110x1110x110x0 : tail0=1'b0;
        16'b10x0x11110x110x0 : tail0=1'b0;
        16'b0x10x11110x110x0 : tail0=1'b0;
        16'b1110x11110x110x0 : tail0=1'b0;
        16'b0x0x111110x110x0 : tail0=1'b0;
        16'b110x111110x110x0 : tail0=1'b0;
        16'b10x1111110x110x0 : tail0=1'b0;
        16'b0x11111110x110x0 : tail0=1'b0;
        16'b1111111110x110x0 : tail0=1'b0;
        16'b0x0x0x0x0x1110x0 : tail0=1'b0;
        16'b110x0x0x0x1110x0 : tail0=1'b0;
        16'b10x10x0x0x1110x0 : tail0=1'b0;
        16'b0x110x0x0x1110x0 : tail0=1'b0;
        16'b11110x0x0x1110x0 : tail0=1'b0;
        16'b10x0x10x0x1110x0 : tail0=1'b0;
        16'b0x10x10x0x1110x0 : tail0=1'b0;
        16'b1110x10x0x1110x0 : tail0=1'b0;
        16'b0x0x110x0x1110x0 : tail0=1'b0;
        16'b110x110x0x1110x0 : tail0=1'b0;
        16'b10x1110x0x1110x0 : tail0=1'b0;
        16'b0x11110x0x1110x0 : tail0=1'b0;
        16'b1111110x0x1110x0 : tail0=1'b0;
        16'b10x0x0x10x1110x0 : tail0=1'b0;
        16'b0x10x0x10x1110x0 : tail0=1'b0;
        16'b1110x0x10x1110x0 : tail0=1'b0;
        16'b0x0x10x10x1110x0 : tail0=1'b0;
        16'b110x10x10x1110x0 : tail0=1'b0;
        16'b10x110x10x1110x0 : tail0=1'b0;
        16'b0x1110x10x1110x0 : tail0=1'b0;
        16'b111110x10x1110x0 : tail0=1'b0;
        16'b0x0x0x110x1110x0 : tail0=1'b0;
        16'b110x0x110x1110x0 : tail0=1'b0;
        16'b10x10x110x1110x0 : tail0=1'b0;
        16'b0x110x110x1110x0 : tail0=1'b0;
        16'b11110x110x1110x0 : tail0=1'b0;
        16'b10x0x1110x1110x0 : tail0=1'b0;
        16'b0x10x1110x1110x0 : tail0=1'b0;
        16'b1110x1110x1110x0 : tail0=1'b0;
        16'b0x0x11110x1110x0 : tail0=1'b0;
        16'b110x11110x1110x0 : tail0=1'b0;
        16'b10x111110x1110x0 : tail0=1'b0;
        16'b0x1111110x1110x0 : tail0=1'b0;
        16'b111111110x1110x0 : tail0=1'b0;
        16'b10x0x0x0x11110x0 : tail0=1'b0;
        16'b0x10x0x0x11110x0 : tail0=1'b0;
        16'b1110x0x0x11110x0 : tail0=1'b0;
        16'b0x0x10x0x11110x0 : tail0=1'b0;
        16'b110x10x0x11110x0 : tail0=1'b0;
        16'b10x110x0x11110x0 : tail0=1'b0;
        16'b0x1110x0x11110x0 : tail0=1'b0;
        16'b111110x0x11110x0 : tail0=1'b0;
        16'b0x0x0x10x11110x0 : tail0=1'b0;
        16'b110x0x10x11110x0 : tail0=1'b0;
        16'b10x10x10x11110x0 : tail0=1'b0;
        16'b0x110x10x11110x0 : tail0=1'b0;
        16'b11110x10x11110x0 : tail0=1'b0;
        16'b10x0x110x11110x0 : tail0=1'b0;
        16'b0x10x110x11110x0 : tail0=1'b0;
        16'b1110x110x11110x0 : tail0=1'b0;
        16'b0x0x1110x11110x0 : tail0=1'b0;
        16'b110x1110x11110x0 : tail0=1'b0;
        16'b10x11110x11110x0 : tail0=1'b0;
        16'b0x111110x11110x0 : tail0=1'b0;
        16'b11111110x11110x0 : tail0=1'b0;
        16'b0x0x0x0x111110x0 : tail0=1'b0;
        16'b110x0x0x111110x0 : tail0=1'b0;
        16'b10x10x0x111110x0 : tail0=1'b0;
        16'b0x110x0x111110x0 : tail0=1'b0;
        16'b11110x0x111110x0 : tail0=1'b0;
        16'b10x0x10x111110x0 : tail0=1'b0;
        16'b0x10x10x111110x0 : tail0=1'b0;
        16'b1110x10x111110x0 : tail0=1'b0;
        16'b0x0x110x111110x0 : tail0=1'b0;
        16'b110x110x111110x0 : tail0=1'b0;
        16'b10x1110x111110x0 : tail0=1'b0;
        16'b0x11110x111110x0 : tail0=1'b0;
        16'b1111110x111110x0 : tail0=1'b0;
        16'b10x0x0x1111110x0 : tail0=1'b0;
        16'b0x10x0x1111110x0 : tail0=1'b0;
        16'b1110x0x1111110x0 : tail0=1'b0;
        16'b0x0x10x1111110x0 : tail0=1'b0;
        16'b110x10x1111110x0 : tail0=1'b0;
        16'b10x110x1111110x0 : tail0=1'b0;
        16'b0x1110x1111110x0 : tail0=1'b0;
        16'b111110x1111110x0 : tail0=1'b0;
        16'b0x0x0x11111110x0 : tail0=1'b0;
        16'b110x0x11111110x0 : tail0=1'b0;
        16'b10x10x11111110x0 : tail0=1'b0;
        16'b0x110x11111110x0 : tail0=1'b0;
        16'b11110x11111110x0 : tail0=1'b0;
        16'b10x0x111111110x0 : tail0=1'b0;
        16'b0x10x111111110x0 : tail0=1'b0;
        16'b1110x111111110x0 : tail0=1'b0;
        16'b0x0x1111111110x0 : tail0=1'b0;
        16'b110x1111111110x0 : tail0=1'b0;
        16'b10x11111111110x0 : tail0=1'b0;
        16'b0x111111111110x0 : tail0=1'b0;
        16'b11111111111110x0 : tail0=1'b0;
        16'b10x0x0x0x0x0x10x : tail0=1'b0;
        16'b0x10x0x0x0x0x10x : tail0=1'b0;
        16'b1110x0x0x0x0x10x : tail0=1'b0;
        16'b0x0x10x0x0x0x10x : tail0=1'b0;
        16'b110x10x0x0x0x10x : tail0=1'b0;
        16'b10x110x0x0x0x10x : tail0=1'b0;
        16'b0x1110x0x0x0x10x : tail0=1'b0;
        16'b111110x0x0x0x10x : tail0=1'b0;
        16'b0x0x0x10x0x0x10x : tail0=1'b0;
        16'b110x0x10x0x0x10x : tail0=1'b0;
        16'b10x10x10x0x0x10x : tail0=1'b0;
        16'b0x110x10x0x0x10x : tail0=1'b0;
        16'b11110x10x0x0x10x : tail0=1'b0;
        16'b10x0x110x0x0x10x : tail0=1'b0;
        16'b0x10x110x0x0x10x : tail0=1'b0;
        16'b1110x110x0x0x10x : tail0=1'b0;
        16'b0x0x1110x0x0x10x : tail0=1'b0;
        16'b110x1110x0x0x10x : tail0=1'b0;
        16'b10x11110x0x0x10x : tail0=1'b0;
        16'b0x111110x0x0x10x : tail0=1'b0;
        16'b11111110x0x0x10x : tail0=1'b0;
        16'b0x0x0x0x10x0x10x : tail0=1'b0;
        16'b110x0x0x10x0x10x : tail0=1'b0;
        16'b10x10x0x10x0x10x : tail0=1'b0;
        16'b0x110x0x10x0x10x : tail0=1'b0;
        16'b11110x0x10x0x10x : tail0=1'b0;
        16'b10x0x10x10x0x10x : tail0=1'b0;
        16'b0x10x10x10x0x10x : tail0=1'b0;
        16'b1110x10x10x0x10x : tail0=1'b0;
        16'b0x0x110x10x0x10x : tail0=1'b0;
        16'b110x110x10x0x10x : tail0=1'b0;
        16'b10x1110x10x0x10x : tail0=1'b0;
        16'b0x11110x10x0x10x : tail0=1'b0;
        16'b1111110x10x0x10x : tail0=1'b0;
        16'b10x0x0x110x0x10x : tail0=1'b0;
        16'b0x10x0x110x0x10x : tail0=1'b0;
        16'b1110x0x110x0x10x : tail0=1'b0;
        16'b0x0x10x110x0x10x : tail0=1'b0;
        16'b110x10x110x0x10x : tail0=1'b0;
        16'b10x110x110x0x10x : tail0=1'b0;
        16'b0x1110x110x0x10x : tail0=1'b0;
        16'b111110x110x0x10x : tail0=1'b0;
        16'b0x0x0x1110x0x10x : tail0=1'b0;
        16'b110x0x1110x0x10x : tail0=1'b0;
        16'b10x10x1110x0x10x : tail0=1'b0;
        16'b0x110x1110x0x10x : tail0=1'b0;
        16'b11110x1110x0x10x : tail0=1'b0;
        16'b10x0x11110x0x10x : tail0=1'b0;
        16'b0x10x11110x0x10x : tail0=1'b0;
        16'b1110x11110x0x10x : tail0=1'b0;
        16'b0x0x111110x0x10x : tail0=1'b0;
        16'b110x111110x0x10x : tail0=1'b0;
        16'b10x1111110x0x10x : tail0=1'b0;
        16'b0x11111110x0x10x : tail0=1'b0;
        16'b1111111110x0x10x : tail0=1'b0;
        16'b0x0x0x0x0x10x10x : tail0=1'b0;
        16'b110x0x0x0x10x10x : tail0=1'b0;
        16'b10x10x0x0x10x10x : tail0=1'b0;
        16'b0x110x0x0x10x10x : tail0=1'b0;
        16'b11110x0x0x10x10x : tail0=1'b0;
        16'b10x0x10x0x10x10x : tail0=1'b0;
        16'b0x10x10x0x10x10x : tail0=1'b0;
        16'b1110x10x0x10x10x : tail0=1'b0;
        16'b0x0x110x0x10x10x : tail0=1'b0;
        16'b110x110x0x10x10x : tail0=1'b0;
        16'b10x1110x0x10x10x : tail0=1'b0;
        16'b0x11110x0x10x10x : tail0=1'b0;
        16'b1111110x0x10x10x : tail0=1'b0;
        16'b10x0x0x10x10x10x : tail0=1'b0;
        16'b0x10x0x10x10x10x : tail0=1'b0;
        16'b1110x0x10x10x10x : tail0=1'b0;
        16'b0x0x10x10x10x10x : tail0=1'b0;
        16'b110x10x10x10x10x : tail0=1'b0;
        16'b10x110x10x10x10x : tail0=1'b0;
        16'b0x1110x10x10x10x : tail0=1'b0;
        16'b111110x10x10x10x : tail0=1'b0;
        16'b0x0x0x110x10x10x : tail0=1'b0;
        16'b110x0x110x10x10x : tail0=1'b0;
        16'b10x10x110x10x10x : tail0=1'b0;
        16'b0x110x110x10x10x : tail0=1'b0;
        16'b11110x110x10x10x : tail0=1'b0;
        16'b10x0x1110x10x10x : tail0=1'b0;
        16'b0x10x1110x10x10x : tail0=1'b0;
        16'b1110x1110x10x10x : tail0=1'b0;
        16'b0x0x11110x10x10x : tail0=1'b0;
        16'b110x11110x10x10x : tail0=1'b0;
        16'b10x111110x10x10x : tail0=1'b0;
        16'b0x1111110x10x10x : tail0=1'b0;
        16'b111111110x10x10x : tail0=1'b0;
        16'b10x0x0x0x110x10x : tail0=1'b0;
        16'b0x10x0x0x110x10x : tail0=1'b0;
        16'b1110x0x0x110x10x : tail0=1'b0;
        16'b0x0x10x0x110x10x : tail0=1'b0;
        16'b110x10x0x110x10x : tail0=1'b0;
        16'b10x110x0x110x10x : tail0=1'b0;
        16'b0x1110x0x110x10x : tail0=1'b0;
        16'b111110x0x110x10x : tail0=1'b0;
        16'b0x0x0x10x110x10x : tail0=1'b0;
        16'b110x0x10x110x10x : tail0=1'b0;
        16'b10x10x10x110x10x : tail0=1'b0;
        16'b0x110x10x110x10x : tail0=1'b0;
        16'b11110x10x110x10x : tail0=1'b0;
        16'b10x0x110x110x10x : tail0=1'b0;
        16'b0x10x110x110x10x : tail0=1'b0;
        16'b1110x110x110x10x : tail0=1'b0;
        16'b0x0x1110x110x10x : tail0=1'b0;
        16'b110x1110x110x10x : tail0=1'b0;
        16'b10x11110x110x10x : tail0=1'b0;
        16'b0x111110x110x10x : tail0=1'b0;
        16'b11111110x110x10x : tail0=1'b0;
        16'b0x0x0x0x1110x10x : tail0=1'b0;
        16'b110x0x0x1110x10x : tail0=1'b0;
        16'b10x10x0x1110x10x : tail0=1'b0;
        16'b0x110x0x1110x10x : tail0=1'b0;
        16'b11110x0x1110x10x : tail0=1'b0;
        16'b10x0x10x1110x10x : tail0=1'b0;
        16'b0x10x10x1110x10x : tail0=1'b0;
        16'b1110x10x1110x10x : tail0=1'b0;
        16'b0x0x110x1110x10x : tail0=1'b0;
        16'b110x110x1110x10x : tail0=1'b0;
        16'b10x1110x1110x10x : tail0=1'b0;
        16'b0x11110x1110x10x : tail0=1'b0;
        16'b1111110x1110x10x : tail0=1'b0;
        16'b10x0x0x11110x10x : tail0=1'b0;
        16'b0x10x0x11110x10x : tail0=1'b0;
        16'b1110x0x11110x10x : tail0=1'b0;
        16'b0x0x10x11110x10x : tail0=1'b0;
        16'b110x10x11110x10x : tail0=1'b0;
        16'b10x110x11110x10x : tail0=1'b0;
        16'b0x1110x11110x10x : tail0=1'b0;
        16'b111110x11110x10x : tail0=1'b0;
        16'b0x0x0x111110x10x : tail0=1'b0;
        16'b110x0x111110x10x : tail0=1'b0;
        16'b10x10x111110x10x : tail0=1'b0;
        16'b0x110x111110x10x : tail0=1'b0;
        16'b11110x111110x10x : tail0=1'b0;
        16'b10x0x1111110x10x : tail0=1'b0;
        16'b0x10x1111110x10x : tail0=1'b0;
        16'b1110x1111110x10x : tail0=1'b0;
        16'b0x0x11111110x10x : tail0=1'b0;
        16'b110x11111110x10x : tail0=1'b0;
        16'b10x111111110x10x : tail0=1'b0;
        16'b0x1111111110x10x : tail0=1'b0;
        16'b111111111110x10x : tail0=1'b0;
        16'b0x0x0x0x0x0x110x : tail0=1'b0;
        16'b110x0x0x0x0x110x : tail0=1'b0;
        16'b10x10x0x0x0x110x : tail0=1'b0;
        16'b0x110x0x0x0x110x : tail0=1'b0;
        16'b11110x0x0x0x110x : tail0=1'b0;
        16'b10x0x10x0x0x110x : tail0=1'b0;
        16'b0x10x10x0x0x110x : tail0=1'b0;
        16'b1110x10x0x0x110x : tail0=1'b0;
        16'b0x0x110x0x0x110x : tail0=1'b0;
        16'b110x110x0x0x110x : tail0=1'b0;
        16'b10x1110x0x0x110x : tail0=1'b0;
        16'b0x11110x0x0x110x : tail0=1'b0;
        16'b1111110x0x0x110x : tail0=1'b0;
        16'b10x0x0x10x0x110x : tail0=1'b0;
        16'b0x10x0x10x0x110x : tail0=1'b0;
        16'b1110x0x10x0x110x : tail0=1'b0;
        16'b0x0x10x10x0x110x : tail0=1'b0;
        16'b110x10x10x0x110x : tail0=1'b0;
        16'b10x110x10x0x110x : tail0=1'b0;
        16'b0x1110x10x0x110x : tail0=1'b0;
        16'b111110x10x0x110x : tail0=1'b0;
        16'b0x0x0x110x0x110x : tail0=1'b0;
        16'b110x0x110x0x110x : tail0=1'b0;
        16'b10x10x110x0x110x : tail0=1'b0;
        16'b0x110x110x0x110x : tail0=1'b0;
        16'b11110x110x0x110x : tail0=1'b0;
        16'b10x0x1110x0x110x : tail0=1'b0;
        16'b0x10x1110x0x110x : tail0=1'b0;
        16'b1110x1110x0x110x : tail0=1'b0;
        16'b0x0x11110x0x110x : tail0=1'b0;
        16'b110x11110x0x110x : tail0=1'b0;
        16'b10x111110x0x110x : tail0=1'b0;
        16'b0x1111110x0x110x : tail0=1'b0;
        16'b111111110x0x110x : tail0=1'b0;
        16'b10x0x0x0x10x110x : tail0=1'b0;
        16'b0x10x0x0x10x110x : tail0=1'b0;
        16'b1110x0x0x10x110x : tail0=1'b0;
        16'b0x0x10x0x10x110x : tail0=1'b0;
        16'b110x10x0x10x110x : tail0=1'b0;
        16'b10x110x0x10x110x : tail0=1'b0;
        16'b0x1110x0x10x110x : tail0=1'b0;
        16'b111110x0x10x110x : tail0=1'b0;
        16'b0x0x0x10x10x110x : tail0=1'b0;
        16'b110x0x10x10x110x : tail0=1'b0;
        16'b10x10x10x10x110x : tail0=1'b0;
        16'b0x110x10x10x110x : tail0=1'b0;
        16'b11110x10x10x110x : tail0=1'b0;
        16'b10x0x110x10x110x : tail0=1'b0;
        16'b0x10x110x10x110x : tail0=1'b0;
        16'b1110x110x10x110x : tail0=1'b0;
        16'b0x0x1110x10x110x : tail0=1'b0;
        16'b110x1110x10x110x : tail0=1'b0;
        16'b10x11110x10x110x : tail0=1'b0;
        16'b0x111110x10x110x : tail0=1'b0;
        16'b11111110x10x110x : tail0=1'b0;
        16'b0x0x0x0x110x110x : tail0=1'b0;
        16'b110x0x0x110x110x : tail0=1'b0;
        16'b10x10x0x110x110x : tail0=1'b0;
        16'b0x110x0x110x110x : tail0=1'b0;
        16'b11110x0x110x110x : tail0=1'b0;
        16'b10x0x10x110x110x : tail0=1'b0;
        16'b0x10x10x110x110x : tail0=1'b0;
        16'b1110x10x110x110x : tail0=1'b0;
        16'b0x0x110x110x110x : tail0=1'b0;
        16'b110x110x110x110x : tail0=1'b0;
        16'b10x1110x110x110x : tail0=1'b0;
        16'b0x11110x110x110x : tail0=1'b0;
        16'b1111110x110x110x : tail0=1'b0;
        16'b10x0x0x1110x110x : tail0=1'b0;
        16'b0x10x0x1110x110x : tail0=1'b0;
        16'b1110x0x1110x110x : tail0=1'b0;
        16'b0x0x10x1110x110x : tail0=1'b0;
        16'b110x10x1110x110x : tail0=1'b0;
        16'b10x110x1110x110x : tail0=1'b0;
        16'b0x1110x1110x110x : tail0=1'b0;
        16'b111110x1110x110x : tail0=1'b0;
        16'b0x0x0x11110x110x : tail0=1'b0;
        16'b110x0x11110x110x : tail0=1'b0;
        16'b10x10x11110x110x : tail0=1'b0;
        16'b0x110x11110x110x : tail0=1'b0;
        16'b11110x11110x110x : tail0=1'b0;
        16'b10x0x111110x110x : tail0=1'b0;
        16'b0x10x111110x110x : tail0=1'b0;
        16'b1110x111110x110x : tail0=1'b0;
        16'b0x0x1111110x110x : tail0=1'b0;
        16'b110x1111110x110x : tail0=1'b0;
        16'b10x11111110x110x : tail0=1'b0;
        16'b0x111111110x110x : tail0=1'b0;
        16'b11111111110x110x : tail0=1'b0;
        16'b10x0x0x0x0x1110x : tail0=1'b0;
        16'b0x10x0x0x0x1110x : tail0=1'b0;
        16'b1110x0x0x0x1110x : tail0=1'b0;
        16'b0x0x10x0x0x1110x : tail0=1'b0;
        16'b110x10x0x0x1110x : tail0=1'b0;
        16'b10x110x0x0x1110x : tail0=1'b0;
        16'b0x1110x0x0x1110x : tail0=1'b0;
        16'b111110x0x0x1110x : tail0=1'b0;
        16'b0x0x0x10x0x1110x : tail0=1'b0;
        16'b110x0x10x0x1110x : tail0=1'b0;
        16'b10x10x10x0x1110x : tail0=1'b0;
        16'b0x110x10x0x1110x : tail0=1'b0;
        16'b11110x10x0x1110x : tail0=1'b0;
        16'b10x0x110x0x1110x : tail0=1'b0;
        16'b0x10x110x0x1110x : tail0=1'b0;
        16'b1110x110x0x1110x : tail0=1'b0;
        16'b0x0x1110x0x1110x : tail0=1'b0;
        16'b110x1110x0x1110x : tail0=1'b0;
        16'b10x11110x0x1110x : tail0=1'b0;
        16'b0x111110x0x1110x : tail0=1'b0;
        16'b11111110x0x1110x : tail0=1'b0;
        16'b0x0x0x0x10x1110x : tail0=1'b0;
        16'b110x0x0x10x1110x : tail0=1'b0;
        16'b10x10x0x10x1110x : tail0=1'b0;
        16'b0x110x0x10x1110x : tail0=1'b0;
        16'b11110x0x10x1110x : tail0=1'b0;
        16'b10x0x10x10x1110x : tail0=1'b0;
        16'b0x10x10x10x1110x : tail0=1'b0;
        16'b1110x10x10x1110x : tail0=1'b0;
        16'b0x0x110x10x1110x : tail0=1'b0;
        16'b110x110x10x1110x : tail0=1'b0;
        16'b10x1110x10x1110x : tail0=1'b0;
        16'b0x11110x10x1110x : tail0=1'b0;
        16'b1111110x10x1110x : tail0=1'b0;
        16'b10x0x0x110x1110x : tail0=1'b0;
        16'b0x10x0x110x1110x : tail0=1'b0;
        16'b1110x0x110x1110x : tail0=1'b0;
        16'b0x0x10x110x1110x : tail0=1'b0;
        16'b110x10x110x1110x : tail0=1'b0;
        16'b10x110x110x1110x : tail0=1'b0;
        16'b0x1110x110x1110x : tail0=1'b0;
        16'b111110x110x1110x : tail0=1'b0;
        16'b0x0x0x1110x1110x : tail0=1'b0;
        16'b110x0x1110x1110x : tail0=1'b0;
        16'b10x10x1110x1110x : tail0=1'b0;
        16'b0x110x1110x1110x : tail0=1'b0;
        16'b11110x1110x1110x : tail0=1'b0;
        16'b10x0x11110x1110x : tail0=1'b0;
        16'b0x10x11110x1110x : tail0=1'b0;
        16'b1110x11110x1110x : tail0=1'b0;
        16'b0x0x111110x1110x : tail0=1'b0;
        16'b110x111110x1110x : tail0=1'b0;
        16'b10x1111110x1110x : tail0=1'b0;
        16'b0x11111110x1110x : tail0=1'b0;
        16'b1111111110x1110x : tail0=1'b0;
        16'b0x0x0x0x0x11110x : tail0=1'b0;
        16'b110x0x0x0x11110x : tail0=1'b0;
        16'b10x10x0x0x11110x : tail0=1'b0;
        16'b0x110x0x0x11110x : tail0=1'b0;
        16'b11110x0x0x11110x : tail0=1'b0;
        16'b10x0x10x0x11110x : tail0=1'b0;
        16'b0x10x10x0x11110x : tail0=1'b0;
        16'b1110x10x0x11110x : tail0=1'b0;
        16'b0x0x110x0x11110x : tail0=1'b0;
        16'b110x110x0x11110x : tail0=1'b0;
        16'b10x1110x0x11110x : tail0=1'b0;
        16'b0x11110x0x11110x : tail0=1'b0;
        16'b1111110x0x11110x : tail0=1'b0;
        16'b10x0x0x10x11110x : tail0=1'b0;
        16'b0x10x0x10x11110x : tail0=1'b0;
        16'b1110x0x10x11110x : tail0=1'b0;
        16'b0x0x10x10x11110x : tail0=1'b0;
        16'b110x10x10x11110x : tail0=1'b0;
        16'b10x110x10x11110x : tail0=1'b0;
        16'b0x1110x10x11110x : tail0=1'b0;
        16'b111110x10x11110x : tail0=1'b0;
        16'b0x0x0x110x11110x : tail0=1'b0;
        16'b110x0x110x11110x : tail0=1'b0;
        16'b10x10x110x11110x : tail0=1'b0;
        16'b0x110x110x11110x : tail0=1'b0;
        16'b11110x110x11110x : tail0=1'b0;
        16'b10x0x1110x11110x : tail0=1'b0;
        16'b0x10x1110x11110x : tail0=1'b0;
        16'b1110x1110x11110x : tail0=1'b0;
        16'b0x0x11110x11110x : tail0=1'b0;
        16'b110x11110x11110x : tail0=1'b0;
        16'b10x111110x11110x : tail0=1'b0;
        16'b0x1111110x11110x : tail0=1'b0;
        16'b111111110x11110x : tail0=1'b0;
        16'b10x0x0x0x111110x : tail0=1'b0;
        16'b0x10x0x0x111110x : tail0=1'b0;
        16'b1110x0x0x111110x : tail0=1'b0;
        16'b0x0x10x0x111110x : tail0=1'b0;
        16'b110x10x0x111110x : tail0=1'b0;
        16'b10x110x0x111110x : tail0=1'b0;
        16'b0x1110x0x111110x : tail0=1'b0;
        16'b111110x0x111110x : tail0=1'b0;
        16'b0x0x0x10x111110x : tail0=1'b0;
        16'b110x0x10x111110x : tail0=1'b0;
        16'b10x10x10x111110x : tail0=1'b0;
        16'b0x110x10x111110x : tail0=1'b0;
        16'b11110x10x111110x : tail0=1'b0;
        16'b10x0x110x111110x : tail0=1'b0;
        16'b0x10x110x111110x : tail0=1'b0;
        16'b1110x110x111110x : tail0=1'b0;
        16'b0x0x1110x111110x : tail0=1'b0;
        16'b110x1110x111110x : tail0=1'b0;
        16'b10x11110x111110x : tail0=1'b0;
        16'b0x111110x111110x : tail0=1'b0;
        16'b11111110x111110x : tail0=1'b0;
        16'b0x0x0x0x1111110x : tail0=1'b0;
        16'b110x0x0x1111110x : tail0=1'b0;
        16'b10x10x0x1111110x : tail0=1'b0;
        16'b0x110x0x1111110x : tail0=1'b0;
        16'b11110x0x1111110x : tail0=1'b0;
        16'b10x0x10x1111110x : tail0=1'b0;
        16'b0x10x10x1111110x : tail0=1'b0;
        16'b1110x10x1111110x : tail0=1'b0;
        16'b0x0x110x1111110x : tail0=1'b0;
        16'b110x110x1111110x : tail0=1'b0;
        16'b10x1110x1111110x : tail0=1'b0;
        16'b0x11110x1111110x : tail0=1'b0;
        16'b1111110x1111110x : tail0=1'b0;
        16'b10x0x0x11111110x : tail0=1'b0;
        16'b0x10x0x11111110x : tail0=1'b0;
        16'b1110x0x11111110x : tail0=1'b0;
        16'b0x0x10x11111110x : tail0=1'b0;
        16'b110x10x11111110x : tail0=1'b0;
        16'b10x110x11111110x : tail0=1'b0;
        16'b0x1110x11111110x : tail0=1'b0;
        16'b111110x11111110x : tail0=1'b0;
        16'b0x0x0x111111110x : tail0=1'b0;
        16'b110x0x111111110x : tail0=1'b0;
        16'b10x10x111111110x : tail0=1'b0;
        16'b0x110x111111110x : tail0=1'b0;
        16'b11110x111111110x : tail0=1'b0;
        16'b10x0x1111111110x : tail0=1'b0;
        16'b0x10x1111111110x : tail0=1'b0;
        16'b1110x1111111110x : tail0=1'b0;
        16'b0x0x11111111110x : tail0=1'b0;
        16'b110x11111111110x : tail0=1'b0;
        16'b10x111111111110x : tail0=1'b0;
        16'b0x1111111111110x : tail0=1'b0;
        16'b111111111111110x : tail0=1'b0;
        16'b0x0x0x0x0x0x0x10 : tail0=1'b0;
        16'b110x0x0x0x0x0x10 : tail0=1'b0;
        16'b10x10x0x0x0x0x10 : tail0=1'b0;
        16'b0x110x0x0x0x0x10 : tail0=1'b0;
        16'b11110x0x0x0x0x10 : tail0=1'b0;
        16'b10x0x10x0x0x0x10 : tail0=1'b0;
        16'b0x10x10x0x0x0x10 : tail0=1'b0;
        16'b1110x10x0x0x0x10 : tail0=1'b0;
        16'b0x0x110x0x0x0x10 : tail0=1'b0;
        16'b110x110x0x0x0x10 : tail0=1'b0;
        16'b10x1110x0x0x0x10 : tail0=1'b0;
        16'b0x11110x0x0x0x10 : tail0=1'b0;
        16'b1111110x0x0x0x10 : tail0=1'b0;
        16'b10x0x0x10x0x0x10 : tail0=1'b0;
        16'b0x10x0x10x0x0x10 : tail0=1'b0;
        16'b1110x0x10x0x0x10 : tail0=1'b0;
        16'b0x0x10x10x0x0x10 : tail0=1'b0;
        16'b110x10x10x0x0x10 : tail0=1'b0;
        16'b10x110x10x0x0x10 : tail0=1'b0;
        16'b0x1110x10x0x0x10 : tail0=1'b0;
        16'b111110x10x0x0x10 : tail0=1'b0;
        16'b0x0x0x110x0x0x10 : tail0=1'b0;
        16'b110x0x110x0x0x10 : tail0=1'b0;
        16'b10x10x110x0x0x10 : tail0=1'b0;
        16'b0x110x110x0x0x10 : tail0=1'b0;
        16'b11110x110x0x0x10 : tail0=1'b0;
        16'b10x0x1110x0x0x10 : tail0=1'b0;
        16'b0x10x1110x0x0x10 : tail0=1'b0;
        16'b1110x1110x0x0x10 : tail0=1'b0;
        16'b0x0x11110x0x0x10 : tail0=1'b0;
        16'b110x11110x0x0x10 : tail0=1'b0;
        16'b10x111110x0x0x10 : tail0=1'b0;
        16'b0x1111110x0x0x10 : tail0=1'b0;
        16'b111111110x0x0x10 : tail0=1'b0;
        16'b10x0x0x0x10x0x10 : tail0=1'b0;
        16'b0x10x0x0x10x0x10 : tail0=1'b0;
        16'b1110x0x0x10x0x10 : tail0=1'b0;
        16'b0x0x10x0x10x0x10 : tail0=1'b0;
        16'b110x10x0x10x0x10 : tail0=1'b0;
        16'b10x110x0x10x0x10 : tail0=1'b0;
        16'b0x1110x0x10x0x10 : tail0=1'b0;
        16'b111110x0x10x0x10 : tail0=1'b0;
        16'b0x0x0x10x10x0x10 : tail0=1'b0;
        16'b110x0x10x10x0x10 : tail0=1'b0;
        16'b10x10x10x10x0x10 : tail0=1'b0;
        16'b0x110x10x10x0x10 : tail0=1'b0;
        16'b11110x10x10x0x10 : tail0=1'b0;
        16'b10x0x110x10x0x10 : tail0=1'b0;
        16'b0x10x110x10x0x10 : tail0=1'b0;
        16'b1110x110x10x0x10 : tail0=1'b0;
        16'b0x0x1110x10x0x10 : tail0=1'b0;
        16'b110x1110x10x0x10 : tail0=1'b0;
        16'b10x11110x10x0x10 : tail0=1'b0;
        16'b0x111110x10x0x10 : tail0=1'b0;
        16'b11111110x10x0x10 : tail0=1'b0;
        16'b0x0x0x0x110x0x10 : tail0=1'b0;
        16'b110x0x0x110x0x10 : tail0=1'b0;
        16'b10x10x0x110x0x10 : tail0=1'b0;
        16'b0x110x0x110x0x10 : tail0=1'b0;
        16'b11110x0x110x0x10 : tail0=1'b0;
        16'b10x0x10x110x0x10 : tail0=1'b0;
        16'b0x10x10x110x0x10 : tail0=1'b0;
        16'b1110x10x110x0x10 : tail0=1'b0;
        16'b0x0x110x110x0x10 : tail0=1'b0;
        16'b110x110x110x0x10 : tail0=1'b0;
        16'b10x1110x110x0x10 : tail0=1'b0;
        16'b0x11110x110x0x10 : tail0=1'b0;
        16'b1111110x110x0x10 : tail0=1'b0;
        16'b10x0x0x1110x0x10 : tail0=1'b0;
        16'b0x10x0x1110x0x10 : tail0=1'b0;
        16'b1110x0x1110x0x10 : tail0=1'b0;
        16'b0x0x10x1110x0x10 : tail0=1'b0;
        16'b110x10x1110x0x10 : tail0=1'b0;
        16'b10x110x1110x0x10 : tail0=1'b0;
        16'b0x1110x1110x0x10 : tail0=1'b0;
        16'b111110x1110x0x10 : tail0=1'b0;
        16'b0x0x0x11110x0x10 : tail0=1'b0;
        16'b110x0x11110x0x10 : tail0=1'b0;
        16'b10x10x11110x0x10 : tail0=1'b0;
        16'b0x110x11110x0x10 : tail0=1'b0;
        16'b11110x11110x0x10 : tail0=1'b0;
        16'b10x0x111110x0x10 : tail0=1'b0;
        16'b0x10x111110x0x10 : tail0=1'b0;
        16'b1110x111110x0x10 : tail0=1'b0;
        16'b0x0x1111110x0x10 : tail0=1'b0;
        16'b110x1111110x0x10 : tail0=1'b0;
        16'b10x11111110x0x10 : tail0=1'b0;
        16'b0x111111110x0x10 : tail0=1'b0;
        16'b11111111110x0x10 : tail0=1'b0;
        16'b10x0x0x0x0x10x10 : tail0=1'b0;
        16'b0x10x0x0x0x10x10 : tail0=1'b0;
        16'b1110x0x0x0x10x10 : tail0=1'b0;
        16'b0x0x10x0x0x10x10 : tail0=1'b0;
        16'b110x10x0x0x10x10 : tail0=1'b0;
        16'b10x110x0x0x10x10 : tail0=1'b0;
        16'b0x1110x0x0x10x10 : tail0=1'b0;
        16'b111110x0x0x10x10 : tail0=1'b0;
        16'b0x0x0x10x0x10x10 : tail0=1'b0;
        16'b110x0x10x0x10x10 : tail0=1'b0;
        16'b10x10x10x0x10x10 : tail0=1'b0;
        16'b0x110x10x0x10x10 : tail0=1'b0;
        16'b11110x10x0x10x10 : tail0=1'b0;
        16'b10x0x110x0x10x10 : tail0=1'b0;
        16'b0x10x110x0x10x10 : tail0=1'b0;
        16'b1110x110x0x10x10 : tail0=1'b0;
        16'b0x0x1110x0x10x10 : tail0=1'b0;
        16'b110x1110x0x10x10 : tail0=1'b0;
        16'b10x11110x0x10x10 : tail0=1'b0;
        16'b0x111110x0x10x10 : tail0=1'b0;
        16'b11111110x0x10x10 : tail0=1'b0;
        16'b0x0x0x0x10x10x10 : tail0=1'b0;
        16'b110x0x0x10x10x10 : tail0=1'b0;
        16'b10x10x0x10x10x10 : tail0=1'b0;
        16'b0x110x0x10x10x10 : tail0=1'b0;
        16'b11110x0x10x10x10 : tail0=1'b0;
        16'b10x0x10x10x10x10 : tail0=1'b0;
        16'b0x10x10x10x10x10 : tail0=1'b0;
        16'b1110x10x10x10x10 : tail0=1'b0;
        16'b0x0x110x10x10x10 : tail0=1'b0;
        16'b110x110x10x10x10 : tail0=1'b0;
        16'b10x1110x10x10x10 : tail0=1'b0;
        16'b0x11110x10x10x10 : tail0=1'b0;
        16'b1111110x10x10x10 : tail0=1'b0;
        16'b10x0x0x110x10x10 : tail0=1'b0;
        16'b0x10x0x110x10x10 : tail0=1'b0;
        16'b1110x0x110x10x10 : tail0=1'b0;
        16'b0x0x10x110x10x10 : tail0=1'b0;
        16'b110x10x110x10x10 : tail0=1'b0;
        16'b10x110x110x10x10 : tail0=1'b0;
        16'b0x1110x110x10x10 : tail0=1'b0;
        16'b111110x110x10x10 : tail0=1'b0;
        16'b0x0x0x1110x10x10 : tail0=1'b0;
        16'b110x0x1110x10x10 : tail0=1'b0;
        16'b10x10x1110x10x10 : tail0=1'b0;
        16'b0x110x1110x10x10 : tail0=1'b0;
        16'b11110x1110x10x10 : tail0=1'b0;
        16'b10x0x11110x10x10 : tail0=1'b0;
        16'b0x10x11110x10x10 : tail0=1'b0;
        16'b1110x11110x10x10 : tail0=1'b0;
        16'b0x0x111110x10x10 : tail0=1'b0;
        16'b110x111110x10x10 : tail0=1'b0;
        16'b10x1111110x10x10 : tail0=1'b0;
        16'b0x11111110x10x10 : tail0=1'b0;
        16'b1111111110x10x10 : tail0=1'b0;
        16'b0x0x0x0x0x110x10 : tail0=1'b0;
        16'b110x0x0x0x110x10 : tail0=1'b0;
        16'b10x10x0x0x110x10 : tail0=1'b0;
        16'b0x110x0x0x110x10 : tail0=1'b0;
        16'b11110x0x0x110x10 : tail0=1'b0;
        16'b10x0x10x0x110x10 : tail0=1'b0;
        16'b0x10x10x0x110x10 : tail0=1'b0;
        16'b1110x10x0x110x10 : tail0=1'b0;
        16'b0x0x110x0x110x10 : tail0=1'b0;
        16'b110x110x0x110x10 : tail0=1'b0;
        16'b10x1110x0x110x10 : tail0=1'b0;
        16'b0x11110x0x110x10 : tail0=1'b0;
        16'b1111110x0x110x10 : tail0=1'b0;
        16'b10x0x0x10x110x10 : tail0=1'b0;
        16'b0x10x0x10x110x10 : tail0=1'b0;
        16'b1110x0x10x110x10 : tail0=1'b0;
        16'b0x0x10x10x110x10 : tail0=1'b0;
        16'b110x10x10x110x10 : tail0=1'b0;
        16'b10x110x10x110x10 : tail0=1'b0;
        16'b0x1110x10x110x10 : tail0=1'b0;
        16'b111110x10x110x10 : tail0=1'b0;
        16'b0x0x0x110x110x10 : tail0=1'b0;
        16'b110x0x110x110x10 : tail0=1'b0;
        16'b10x10x110x110x10 : tail0=1'b0;
        16'b0x110x110x110x10 : tail0=1'b0;
        16'b11110x110x110x10 : tail0=1'b0;
        16'b10x0x1110x110x10 : tail0=1'b0;
        16'b0x10x1110x110x10 : tail0=1'b0;
        16'b1110x1110x110x10 : tail0=1'b0;
        16'b0x0x11110x110x10 : tail0=1'b0;
        16'b110x11110x110x10 : tail0=1'b0;
        16'b10x111110x110x10 : tail0=1'b0;
        16'b0x1111110x110x10 : tail0=1'b0;
        16'b111111110x110x10 : tail0=1'b0;
        16'b10x0x0x0x1110x10 : tail0=1'b0;
        16'b0x10x0x0x1110x10 : tail0=1'b0;
        16'b1110x0x0x1110x10 : tail0=1'b0;
        16'b0x0x10x0x1110x10 : tail0=1'b0;
        16'b110x10x0x1110x10 : tail0=1'b0;
        16'b10x110x0x1110x10 : tail0=1'b0;
        16'b0x1110x0x1110x10 : tail0=1'b0;
        16'b111110x0x1110x10 : tail0=1'b0;
        16'b0x0x0x10x1110x10 : tail0=1'b0;
        16'b110x0x10x1110x10 : tail0=1'b0;
        16'b10x10x10x1110x10 : tail0=1'b0;
        16'b0x110x10x1110x10 : tail0=1'b0;
        16'b11110x10x1110x10 : tail0=1'b0;
        16'b10x0x110x1110x10 : tail0=1'b0;
        16'b0x10x110x1110x10 : tail0=1'b0;
        16'b1110x110x1110x10 : tail0=1'b0;
        16'b0x0x1110x1110x10 : tail0=1'b0;
        16'b110x1110x1110x10 : tail0=1'b0;
        16'b10x11110x1110x10 : tail0=1'b0;
        16'b0x111110x1110x10 : tail0=1'b0;
        16'b11111110x1110x10 : tail0=1'b0;
        16'b0x0x0x0x11110x10 : tail0=1'b0;
        16'b110x0x0x11110x10 : tail0=1'b0;
        16'b10x10x0x11110x10 : tail0=1'b0;
        16'b0x110x0x11110x10 : tail0=1'b0;
        16'b11110x0x11110x10 : tail0=1'b0;
        16'b10x0x10x11110x10 : tail0=1'b0;
        16'b0x10x10x11110x10 : tail0=1'b0;
        16'b1110x10x11110x10 : tail0=1'b0;
        16'b0x0x110x11110x10 : tail0=1'b0;
        16'b110x110x11110x10 : tail0=1'b0;
        16'b10x1110x11110x10 : tail0=1'b0;
        16'b0x11110x11110x10 : tail0=1'b0;
        16'b1111110x11110x10 : tail0=1'b0;
        16'b10x0x0x111110x10 : tail0=1'b0;
        16'b0x10x0x111110x10 : tail0=1'b0;
        16'b1110x0x111110x10 : tail0=1'b0;
        16'b0x0x10x111110x10 : tail0=1'b0;
        16'b110x10x111110x10 : tail0=1'b0;
        16'b10x110x111110x10 : tail0=1'b0;
        16'b0x1110x111110x10 : tail0=1'b0;
        16'b111110x111110x10 : tail0=1'b0;
        16'b0x0x0x1111110x10 : tail0=1'b0;
        16'b110x0x1111110x10 : tail0=1'b0;
        16'b10x10x1111110x10 : tail0=1'b0;
        16'b0x110x1111110x10 : tail0=1'b0;
        16'b11110x1111110x10 : tail0=1'b0;
        16'b10x0x11111110x10 : tail0=1'b0;
        16'b0x10x11111110x10 : tail0=1'b0;
        16'b1110x11111110x10 : tail0=1'b0;
        16'b0x0x111111110x10 : tail0=1'b0;
        16'b110x111111110x10 : tail0=1'b0;
        16'b10x1111111110x10 : tail0=1'b0;
        16'b0x11111111110x10 : tail0=1'b0;
        16'b1111111111110x10 : tail0=1'b0;
        16'b10x0x0x0x0x0x110 : tail0=1'b0;
        16'b0x10x0x0x0x0x110 : tail0=1'b0;
        16'b1110x0x0x0x0x110 : tail0=1'b0;
        16'b0x0x10x0x0x0x110 : tail0=1'b0;
        16'b110x10x0x0x0x110 : tail0=1'b0;
        16'b10x110x0x0x0x110 : tail0=1'b0;
        16'b0x1110x0x0x0x110 : tail0=1'b0;
        16'b111110x0x0x0x110 : tail0=1'b0;
        16'b0x0x0x10x0x0x110 : tail0=1'b0;
        16'b110x0x10x0x0x110 : tail0=1'b0;
        16'b10x10x10x0x0x110 : tail0=1'b0;
        16'b0x110x10x0x0x110 : tail0=1'b0;
        16'b11110x10x0x0x110 : tail0=1'b0;
        16'b10x0x110x0x0x110 : tail0=1'b0;
        16'b0x10x110x0x0x110 : tail0=1'b0;
        16'b1110x110x0x0x110 : tail0=1'b0;
        16'b0x0x1110x0x0x110 : tail0=1'b0;
        16'b110x1110x0x0x110 : tail0=1'b0;
        16'b10x11110x0x0x110 : tail0=1'b0;
        16'b0x111110x0x0x110 : tail0=1'b0;
        16'b11111110x0x0x110 : tail0=1'b0;
        16'b0x0x0x0x10x0x110 : tail0=1'b0;
        16'b110x0x0x10x0x110 : tail0=1'b0;
        16'b10x10x0x10x0x110 : tail0=1'b0;
        16'b0x110x0x10x0x110 : tail0=1'b0;
        16'b11110x0x10x0x110 : tail0=1'b0;
        16'b10x0x10x10x0x110 : tail0=1'b0;
        16'b0x10x10x10x0x110 : tail0=1'b0;
        16'b1110x10x10x0x110 : tail0=1'b0;
        16'b0x0x110x10x0x110 : tail0=1'b0;
        16'b110x110x10x0x110 : tail0=1'b0;
        16'b10x1110x10x0x110 : tail0=1'b0;
        16'b0x11110x10x0x110 : tail0=1'b0;
        16'b1111110x10x0x110 : tail0=1'b0;
        16'b10x0x0x110x0x110 : tail0=1'b0;
        16'b0x10x0x110x0x110 : tail0=1'b0;
        16'b1110x0x110x0x110 : tail0=1'b0;
        16'b0x0x10x110x0x110 : tail0=1'b0;
        16'b110x10x110x0x110 : tail0=1'b0;
        16'b10x110x110x0x110 : tail0=1'b0;
        16'b0x1110x110x0x110 : tail0=1'b0;
        16'b111110x110x0x110 : tail0=1'b0;
        16'b0x0x0x1110x0x110 : tail0=1'b0;
        16'b110x0x1110x0x110 : tail0=1'b0;
        16'b10x10x1110x0x110 : tail0=1'b0;
        16'b0x110x1110x0x110 : tail0=1'b0;
        16'b11110x1110x0x110 : tail0=1'b0;
        16'b10x0x11110x0x110 : tail0=1'b0;
        16'b0x10x11110x0x110 : tail0=1'b0;
        16'b1110x11110x0x110 : tail0=1'b0;
        16'b0x0x111110x0x110 : tail0=1'b0;
        16'b110x111110x0x110 : tail0=1'b0;
        16'b10x1111110x0x110 : tail0=1'b0;
        16'b0x11111110x0x110 : tail0=1'b0;
        16'b1111111110x0x110 : tail0=1'b0;
        16'b0x0x0x0x0x10x110 : tail0=1'b0;
        16'b110x0x0x0x10x110 : tail0=1'b0;
        16'b10x10x0x0x10x110 : tail0=1'b0;
        16'b0x110x0x0x10x110 : tail0=1'b0;
        16'b11110x0x0x10x110 : tail0=1'b0;
        16'b10x0x10x0x10x110 : tail0=1'b0;
        16'b0x10x10x0x10x110 : tail0=1'b0;
        16'b1110x10x0x10x110 : tail0=1'b0;
        16'b0x0x110x0x10x110 : tail0=1'b0;
        16'b110x110x0x10x110 : tail0=1'b0;
        16'b10x1110x0x10x110 : tail0=1'b0;
        16'b0x11110x0x10x110 : tail0=1'b0;
        16'b1111110x0x10x110 : tail0=1'b0;
        16'b10x0x0x10x10x110 : tail0=1'b0;
        16'b0x10x0x10x10x110 : tail0=1'b0;
        16'b1110x0x10x10x110 : tail0=1'b0;
        16'b0x0x10x10x10x110 : tail0=1'b0;
        16'b110x10x10x10x110 : tail0=1'b0;
        16'b10x110x10x10x110 : tail0=1'b0;
        16'b0x1110x10x10x110 : tail0=1'b0;
        16'b111110x10x10x110 : tail0=1'b0;
        16'b0x0x0x110x10x110 : tail0=1'b0;
        16'b110x0x110x10x110 : tail0=1'b0;
        16'b10x10x110x10x110 : tail0=1'b0;
        16'b0x110x110x10x110 : tail0=1'b0;
        16'b11110x110x10x110 : tail0=1'b0;
        16'b10x0x1110x10x110 : tail0=1'b0;
        16'b0x10x1110x10x110 : tail0=1'b0;
        16'b1110x1110x10x110 : tail0=1'b0;
        16'b0x0x11110x10x110 : tail0=1'b0;
        16'b110x11110x10x110 : tail0=1'b0;
        16'b10x111110x10x110 : tail0=1'b0;
        16'b0x1111110x10x110 : tail0=1'b0;
        16'b111111110x10x110 : tail0=1'b0;
        16'b10x0x0x0x110x110 : tail0=1'b0;
        16'b0x10x0x0x110x110 : tail0=1'b0;
        16'b1110x0x0x110x110 : tail0=1'b0;
        16'b0x0x10x0x110x110 : tail0=1'b0;
        16'b110x10x0x110x110 : tail0=1'b0;
        16'b10x110x0x110x110 : tail0=1'b0;
        16'b0x1110x0x110x110 : tail0=1'b0;
        16'b111110x0x110x110 : tail0=1'b0;
        16'b0x0x0x10x110x110 : tail0=1'b0;
        16'b110x0x10x110x110 : tail0=1'b0;
        16'b10x10x10x110x110 : tail0=1'b0;
        16'b0x110x10x110x110 : tail0=1'b0;
        16'b11110x10x110x110 : tail0=1'b0;
        16'b10x0x110x110x110 : tail0=1'b0;
        16'b0x10x110x110x110 : tail0=1'b0;
        16'b1110x110x110x110 : tail0=1'b0;
        16'b0x0x1110x110x110 : tail0=1'b0;
        16'b110x1110x110x110 : tail0=1'b0;
        16'b10x11110x110x110 : tail0=1'b0;
        16'b0x111110x110x110 : tail0=1'b0;
        16'b11111110x110x110 : tail0=1'b0;
        16'b0x0x0x0x1110x110 : tail0=1'b0;
        16'b110x0x0x1110x110 : tail0=1'b0;
        16'b10x10x0x1110x110 : tail0=1'b0;
        16'b0x110x0x1110x110 : tail0=1'b0;
        16'b11110x0x1110x110 : tail0=1'b0;
        16'b10x0x10x1110x110 : tail0=1'b0;
        16'b0x10x10x1110x110 : tail0=1'b0;
        16'b1110x10x1110x110 : tail0=1'b0;
        16'b0x0x110x1110x110 : tail0=1'b0;
        16'b110x110x1110x110 : tail0=1'b0;
        16'b10x1110x1110x110 : tail0=1'b0;
        16'b0x11110x1110x110 : tail0=1'b0;
        16'b1111110x1110x110 : tail0=1'b0;
        16'b10x0x0x11110x110 : tail0=1'b0;
        16'b0x10x0x11110x110 : tail0=1'b0;
        16'b1110x0x11110x110 : tail0=1'b0;
        16'b0x0x10x11110x110 : tail0=1'b0;
        16'b110x10x11110x110 : tail0=1'b0;
        16'b10x110x11110x110 : tail0=1'b0;
        16'b0x1110x11110x110 : tail0=1'b0;
        16'b111110x11110x110 : tail0=1'b0;
        16'b0x0x0x111110x110 : tail0=1'b0;
        16'b110x0x111110x110 : tail0=1'b0;
        16'b10x10x111110x110 : tail0=1'b0;
        16'b0x110x111110x110 : tail0=1'b0;
        16'b11110x111110x110 : tail0=1'b0;
        16'b10x0x1111110x110 : tail0=1'b0;
        16'b0x10x1111110x110 : tail0=1'b0;
        16'b1110x1111110x110 : tail0=1'b0;
        16'b0x0x11111110x110 : tail0=1'b0;
        16'b110x11111110x110 : tail0=1'b0;
        16'b10x111111110x110 : tail0=1'b0;
        16'b0x1111111110x110 : tail0=1'b0;
        16'b111111111110x110 : tail0=1'b0;
        16'b0x0x0x0x0x0x1110 : tail0=1'b0;
        16'b110x0x0x0x0x1110 : tail0=1'b0;
        16'b10x10x0x0x0x1110 : tail0=1'b0;
        16'b0x110x0x0x0x1110 : tail0=1'b0;
        16'b11110x0x0x0x1110 : tail0=1'b0;
        16'b10x0x10x0x0x1110 : tail0=1'b0;
        16'b0x10x10x0x0x1110 : tail0=1'b0;
        16'b1110x10x0x0x1110 : tail0=1'b0;
        16'b0x0x110x0x0x1110 : tail0=1'b0;
        16'b110x110x0x0x1110 : tail0=1'b0;
        16'b10x1110x0x0x1110 : tail0=1'b0;
        16'b0x11110x0x0x1110 : tail0=1'b0;
        16'b1111110x0x0x1110 : tail0=1'b0;
        16'b10x0x0x10x0x1110 : tail0=1'b0;
        16'b0x10x0x10x0x1110 : tail0=1'b0;
        16'b1110x0x10x0x1110 : tail0=1'b0;
        16'b0x0x10x10x0x1110 : tail0=1'b0;
        16'b110x10x10x0x1110 : tail0=1'b0;
        16'b10x110x10x0x1110 : tail0=1'b0;
        16'b0x1110x10x0x1110 : tail0=1'b0;
        16'b111110x10x0x1110 : tail0=1'b0;
        16'b0x0x0x110x0x1110 : tail0=1'b0;
        16'b110x0x110x0x1110 : tail0=1'b0;
        16'b10x10x110x0x1110 : tail0=1'b0;
        16'b0x110x110x0x1110 : tail0=1'b0;
        16'b11110x110x0x1110 : tail0=1'b0;
        16'b10x0x1110x0x1110 : tail0=1'b0;
        16'b0x10x1110x0x1110 : tail0=1'b0;
        16'b1110x1110x0x1110 : tail0=1'b0;
        16'b0x0x11110x0x1110 : tail0=1'b0;
        16'b110x11110x0x1110 : tail0=1'b0;
        16'b10x111110x0x1110 : tail0=1'b0;
        16'b0x1111110x0x1110 : tail0=1'b0;
        16'b111111110x0x1110 : tail0=1'b0;
        16'b10x0x0x0x10x1110 : tail0=1'b0;
        16'b0x10x0x0x10x1110 : tail0=1'b0;
        16'b1110x0x0x10x1110 : tail0=1'b0;
        16'b0x0x10x0x10x1110 : tail0=1'b0;
        16'b110x10x0x10x1110 : tail0=1'b0;
        16'b10x110x0x10x1110 : tail0=1'b0;
        16'b0x1110x0x10x1110 : tail0=1'b0;
        16'b111110x0x10x1110 : tail0=1'b0;
        16'b0x0x0x10x10x1110 : tail0=1'b0;
        16'b110x0x10x10x1110 : tail0=1'b0;
        16'b10x10x10x10x1110 : tail0=1'b0;
        16'b0x110x10x10x1110 : tail0=1'b0;
        16'b11110x10x10x1110 : tail0=1'b0;
        16'b10x0x110x10x1110 : tail0=1'b0;
        16'b0x10x110x10x1110 : tail0=1'b0;
        16'b1110x110x10x1110 : tail0=1'b0;
        16'b0x0x1110x10x1110 : tail0=1'b0;
        16'b110x1110x10x1110 : tail0=1'b0;
        16'b10x11110x10x1110 : tail0=1'b0;
        16'b0x111110x10x1110 : tail0=1'b0;
        16'b11111110x10x1110 : tail0=1'b0;
        16'b0x0x0x0x110x1110 : tail0=1'b0;
        16'b110x0x0x110x1110 : tail0=1'b0;
        16'b10x10x0x110x1110 : tail0=1'b0;
        16'b0x110x0x110x1110 : tail0=1'b0;
        16'b11110x0x110x1110 : tail0=1'b0;
        16'b10x0x10x110x1110 : tail0=1'b0;
        16'b0x10x10x110x1110 : tail0=1'b0;
        16'b1110x10x110x1110 : tail0=1'b0;
        16'b0x0x110x110x1110 : tail0=1'b0;
        16'b110x110x110x1110 : tail0=1'b0;
        16'b10x1110x110x1110 : tail0=1'b0;
        16'b0x11110x110x1110 : tail0=1'b0;
        16'b1111110x110x1110 : tail0=1'b0;
        16'b10x0x0x1110x1110 : tail0=1'b0;
        16'b0x10x0x1110x1110 : tail0=1'b0;
        16'b1110x0x1110x1110 : tail0=1'b0;
        16'b0x0x10x1110x1110 : tail0=1'b0;
        16'b110x10x1110x1110 : tail0=1'b0;
        16'b10x110x1110x1110 : tail0=1'b0;
        16'b0x1110x1110x1110 : tail0=1'b0;
        16'b111110x1110x1110 : tail0=1'b0;
        16'b0x0x0x11110x1110 : tail0=1'b0;
        16'b110x0x11110x1110 : tail0=1'b0;
        16'b10x10x11110x1110 : tail0=1'b0;
        16'b0x110x11110x1110 : tail0=1'b0;
        16'b11110x11110x1110 : tail0=1'b0;
        16'b10x0x111110x1110 : tail0=1'b0;
        16'b0x10x111110x1110 : tail0=1'b0;
        16'b1110x111110x1110 : tail0=1'b0;
        16'b0x0x1111110x1110 : tail0=1'b0;
        16'b110x1111110x1110 : tail0=1'b0;
        16'b10x11111110x1110 : tail0=1'b0;
        16'b0x111111110x1110 : tail0=1'b0;
        16'b11111111110x1110 : tail0=1'b0;
        16'b10x0x0x0x0x11110 : tail0=1'b0;
        16'b0x10x0x0x0x11110 : tail0=1'b0;
        16'b1110x0x0x0x11110 : tail0=1'b0;
        16'b0x0x10x0x0x11110 : tail0=1'b0;
        16'b110x10x0x0x11110 : tail0=1'b0;
        16'b10x110x0x0x11110 : tail0=1'b0;
        16'b0x1110x0x0x11110 : tail0=1'b0;
        16'b111110x0x0x11110 : tail0=1'b0;
        16'b0x0x0x10x0x11110 : tail0=1'b0;
        16'b110x0x10x0x11110 : tail0=1'b0;
        16'b10x10x10x0x11110 : tail0=1'b0;
        16'b0x110x10x0x11110 : tail0=1'b0;
        16'b11110x10x0x11110 : tail0=1'b0;
        16'b10x0x110x0x11110 : tail0=1'b0;
        16'b0x10x110x0x11110 : tail0=1'b0;
        16'b1110x110x0x11110 : tail0=1'b0;
        16'b0x0x1110x0x11110 : tail0=1'b0;
        16'b110x1110x0x11110 : tail0=1'b0;
        16'b10x11110x0x11110 : tail0=1'b0;
        16'b0x111110x0x11110 : tail0=1'b0;
        16'b11111110x0x11110 : tail0=1'b0;
        16'b0x0x0x0x10x11110 : tail0=1'b0;
        16'b110x0x0x10x11110 : tail0=1'b0;
        16'b10x10x0x10x11110 : tail0=1'b0;
        16'b0x110x0x10x11110 : tail0=1'b0;
        16'b11110x0x10x11110 : tail0=1'b0;
        16'b10x0x10x10x11110 : tail0=1'b0;
        16'b0x10x10x10x11110 : tail0=1'b0;
        16'b1110x10x10x11110 : tail0=1'b0;
        16'b0x0x110x10x11110 : tail0=1'b0;
        16'b110x110x10x11110 : tail0=1'b0;
        16'b10x1110x10x11110 : tail0=1'b0;
        16'b0x11110x10x11110 : tail0=1'b0;
        16'b1111110x10x11110 : tail0=1'b0;
        16'b10x0x0x110x11110 : tail0=1'b0;
        16'b0x10x0x110x11110 : tail0=1'b0;
        16'b1110x0x110x11110 : tail0=1'b0;
        16'b0x0x10x110x11110 : tail0=1'b0;
        16'b110x10x110x11110 : tail0=1'b0;
        16'b10x110x110x11110 : tail0=1'b0;
        16'b0x1110x110x11110 : tail0=1'b0;
        16'b111110x110x11110 : tail0=1'b0;
        16'b0x0x0x1110x11110 : tail0=1'b0;
        16'b110x0x1110x11110 : tail0=1'b0;
        16'b10x10x1110x11110 : tail0=1'b0;
        16'b0x110x1110x11110 : tail0=1'b0;
        16'b11110x1110x11110 : tail0=1'b0;
        16'b10x0x11110x11110 : tail0=1'b0;
        16'b0x10x11110x11110 : tail0=1'b0;
        16'b1110x11110x11110 : tail0=1'b0;
        16'b0x0x111110x11110 : tail0=1'b0;
        16'b110x111110x11110 : tail0=1'b0;
        16'b10x1111110x11110 : tail0=1'b0;
        16'b0x11111110x11110 : tail0=1'b0;
        16'b1111111110x11110 : tail0=1'b0;
        16'b0x0x0x0x0x111110 : tail0=1'b0;
        16'b110x0x0x0x111110 : tail0=1'b0;
        16'b10x10x0x0x111110 : tail0=1'b0;
        16'b0x110x0x0x111110 : tail0=1'b0;
        16'b11110x0x0x111110 : tail0=1'b0;
        16'b10x0x10x0x111110 : tail0=1'b0;
        16'b0x10x10x0x111110 : tail0=1'b0;
        16'b1110x10x0x111110 : tail0=1'b0;
        16'b0x0x110x0x111110 : tail0=1'b0;
        16'b110x110x0x111110 : tail0=1'b0;
        16'b10x1110x0x111110 : tail0=1'b0;
        16'b0x11110x0x111110 : tail0=1'b0;
        16'b1111110x0x111110 : tail0=1'b0;
        16'b10x0x0x10x111110 : tail0=1'b0;
        16'b0x10x0x10x111110 : tail0=1'b0;
        16'b1110x0x10x111110 : tail0=1'b0;
        16'b0x0x10x10x111110 : tail0=1'b0;
        16'b110x10x10x111110 : tail0=1'b0;
        16'b10x110x10x111110 : tail0=1'b0;
        16'b0x1110x10x111110 : tail0=1'b0;
        16'b111110x10x111110 : tail0=1'b0;
        16'b0x0x0x110x111110 : tail0=1'b0;
        16'b110x0x110x111110 : tail0=1'b0;
        16'b10x10x110x111110 : tail0=1'b0;
        16'b0x110x110x111110 : tail0=1'b0;
        16'b11110x110x111110 : tail0=1'b0;
        16'b10x0x1110x111110 : tail0=1'b0;
        16'b0x10x1110x111110 : tail0=1'b0;
        16'b1110x1110x111110 : tail0=1'b0;
        16'b0x0x11110x111110 : tail0=1'b0;
        16'b110x11110x111110 : tail0=1'b0;
        16'b10x111110x111110 : tail0=1'b0;
        16'b0x1111110x111110 : tail0=1'b0;
        16'b111111110x111110 : tail0=1'b0;
        16'b10x0x0x0x1111110 : tail0=1'b0;
        16'b0x10x0x0x1111110 : tail0=1'b0;
        16'b1110x0x0x1111110 : tail0=1'b0;
        16'b0x0x10x0x1111110 : tail0=1'b0;
        16'b110x10x0x1111110 : tail0=1'b0;
        16'b10x110x0x1111110 : tail0=1'b0;
        16'b0x1110x0x1111110 : tail0=1'b0;
        16'b111110x0x1111110 : tail0=1'b0;
        16'b0x0x0x10x1111110 : tail0=1'b0;
        16'b110x0x10x1111110 : tail0=1'b0;
        16'b10x10x10x1111110 : tail0=1'b0;
        16'b0x110x10x1111110 : tail0=1'b0;
        16'b11110x10x1111110 : tail0=1'b0;
        16'b10x0x110x1111110 : tail0=1'b0;
        16'b0x10x110x1111110 : tail0=1'b0;
        16'b1110x110x1111110 : tail0=1'b0;
        16'b0x0x1110x1111110 : tail0=1'b0;
        16'b110x1110x1111110 : tail0=1'b0;
        16'b10x11110x1111110 : tail0=1'b0;
        16'b0x111110x1111110 : tail0=1'b0;
        16'b11111110x1111110 : tail0=1'b0;
        16'b0x0x0x0x11111110 : tail0=1'b0;
        16'b110x0x0x11111110 : tail0=1'b0;
        16'b10x10x0x11111110 : tail0=1'b0;
        16'b0x110x0x11111110 : tail0=1'b0;
        16'b11110x0x11111110 : tail0=1'b0;
        16'b10x0x10x11111110 : tail0=1'b0;
        16'b0x10x10x11111110 : tail0=1'b0;
        16'b1110x10x11111110 : tail0=1'b0;
        16'b0x0x110x11111110 : tail0=1'b0;
        16'b110x110x11111110 : tail0=1'b0;
        16'b10x1110x11111110 : tail0=1'b0;
        16'b0x11110x11111110 : tail0=1'b0;
        16'b1111110x11111110 : tail0=1'b0;
        16'b10x0x0x111111110 : tail0=1'b0;
        16'b0x10x0x111111110 : tail0=1'b0;
        16'b1110x0x111111110 : tail0=1'b0;
        16'b0x0x10x111111110 : tail0=1'b0;
        16'b110x10x111111110 : tail0=1'b0;
        16'b10x110x111111110 : tail0=1'b0;
        16'b0x1110x111111110 : tail0=1'b0;
        16'b111110x111111110 : tail0=1'b0;
        16'b0x0x0x1111111110 : tail0=1'b0;
        16'b110x0x1111111110 : tail0=1'b0;
        16'b10x10x1111111110 : tail0=1'b0;
        16'b0x110x1111111110 : tail0=1'b0;
        16'b11110x1111111110 : tail0=1'b0;
        16'b10x0x11111111110 : tail0=1'b0;
        16'b0x10x11111111110 : tail0=1'b0;
        16'b1110x11111111110 : tail0=1'b0;
        16'b0x0x111111111110 : tail0=1'b0;
        16'b110x111111111110 : tail0=1'b0;
        16'b10x1111111111110 : tail0=1'b0;
        16'b0x11111111111110 : tail0=1'b0;
        16'b1111111111111110 : tail0=1'b0;
        16'b10x0x0x0x0x0x0x1 : tail0=1'b0;
        16'b0x10x0x0x0x0x0x1 : tail0=1'b0;
        16'b1110x0x0x0x0x0x1 : tail0=1'b0;
        16'b0x0x10x0x0x0x0x1 : tail0=1'b0;
        16'b110x10x0x0x0x0x1 : tail0=1'b0;
        16'b10x110x0x0x0x0x1 : tail0=1'b0;
        16'b0x1110x0x0x0x0x1 : tail0=1'b0;
        16'b111110x0x0x0x0x1 : tail0=1'b0;
        16'b0x0x0x10x0x0x0x1 : tail0=1'b0;
        16'b110x0x10x0x0x0x1 : tail0=1'b0;
        16'b10x10x10x0x0x0x1 : tail0=1'b0;
        16'b0x110x10x0x0x0x1 : tail0=1'b0;
        16'b11110x10x0x0x0x1 : tail0=1'b0;
        16'b10x0x110x0x0x0x1 : tail0=1'b0;
        16'b0x10x110x0x0x0x1 : tail0=1'b0;
        16'b1110x110x0x0x0x1 : tail0=1'b0;
        16'b0x0x1110x0x0x0x1 : tail0=1'b0;
        16'b110x1110x0x0x0x1 : tail0=1'b0;
        16'b10x11110x0x0x0x1 : tail0=1'b0;
        16'b0x111110x0x0x0x1 : tail0=1'b0;
        16'b11111110x0x0x0x1 : tail0=1'b0;
        16'b0x0x0x0x10x0x0x1 : tail0=1'b0;
        16'b110x0x0x10x0x0x1 : tail0=1'b0;
        16'b10x10x0x10x0x0x1 : tail0=1'b0;
        16'b0x110x0x10x0x0x1 : tail0=1'b0;
        16'b11110x0x10x0x0x1 : tail0=1'b0;
        16'b10x0x10x10x0x0x1 : tail0=1'b0;
        16'b0x10x10x10x0x0x1 : tail0=1'b0;
        16'b1110x10x10x0x0x1 : tail0=1'b0;
        16'b0x0x110x10x0x0x1 : tail0=1'b0;
        16'b110x110x10x0x0x1 : tail0=1'b0;
        16'b10x1110x10x0x0x1 : tail0=1'b0;
        16'b0x11110x10x0x0x1 : tail0=1'b0;
        16'b1111110x10x0x0x1 : tail0=1'b0;
        16'b10x0x0x110x0x0x1 : tail0=1'b0;
        16'b0x10x0x110x0x0x1 : tail0=1'b0;
        16'b1110x0x110x0x0x1 : tail0=1'b0;
        16'b0x0x10x110x0x0x1 : tail0=1'b0;
        16'b110x10x110x0x0x1 : tail0=1'b0;
        16'b10x110x110x0x0x1 : tail0=1'b0;
        16'b0x1110x110x0x0x1 : tail0=1'b0;
        16'b111110x110x0x0x1 : tail0=1'b0;
        16'b0x0x0x1110x0x0x1 : tail0=1'b0;
        16'b110x0x1110x0x0x1 : tail0=1'b0;
        16'b10x10x1110x0x0x1 : tail0=1'b0;
        16'b0x110x1110x0x0x1 : tail0=1'b0;
        16'b11110x1110x0x0x1 : tail0=1'b0;
        16'b10x0x11110x0x0x1 : tail0=1'b0;
        16'b0x10x11110x0x0x1 : tail0=1'b0;
        16'b1110x11110x0x0x1 : tail0=1'b0;
        16'b0x0x111110x0x0x1 : tail0=1'b0;
        16'b110x111110x0x0x1 : tail0=1'b0;
        16'b10x1111110x0x0x1 : tail0=1'b0;
        16'b0x11111110x0x0x1 : tail0=1'b0;
        16'b1111111110x0x0x1 : tail0=1'b0;
        16'b0x0x0x0x0x10x0x1 : tail0=1'b0;
        16'b110x0x0x0x10x0x1 : tail0=1'b0;
        16'b10x10x0x0x10x0x1 : tail0=1'b0;
        16'b0x110x0x0x10x0x1 : tail0=1'b0;
        16'b11110x0x0x10x0x1 : tail0=1'b0;
        16'b10x0x10x0x10x0x1 : tail0=1'b0;
        16'b0x10x10x0x10x0x1 : tail0=1'b0;
        16'b1110x10x0x10x0x1 : tail0=1'b0;
        16'b0x0x110x0x10x0x1 : tail0=1'b0;
        16'b110x110x0x10x0x1 : tail0=1'b0;
        16'b10x1110x0x10x0x1 : tail0=1'b0;
        16'b0x11110x0x10x0x1 : tail0=1'b0;
        16'b1111110x0x10x0x1 : tail0=1'b0;
        16'b10x0x0x10x10x0x1 : tail0=1'b0;
        16'b0x10x0x10x10x0x1 : tail0=1'b0;
        16'b1110x0x10x10x0x1 : tail0=1'b0;
        16'b0x0x10x10x10x0x1 : tail0=1'b0;
        16'b110x10x10x10x0x1 : tail0=1'b0;
        16'b10x110x10x10x0x1 : tail0=1'b0;
        16'b0x1110x10x10x0x1 : tail0=1'b0;
        16'b111110x10x10x0x1 : tail0=1'b0;
        16'b0x0x0x110x10x0x1 : tail0=1'b0;
        16'b110x0x110x10x0x1 : tail0=1'b0;
        16'b10x10x110x10x0x1 : tail0=1'b0;
        16'b0x110x110x10x0x1 : tail0=1'b0;
        16'b11110x110x10x0x1 : tail0=1'b0;
        16'b10x0x1110x10x0x1 : tail0=1'b0;
        16'b0x10x1110x10x0x1 : tail0=1'b0;
        16'b1110x1110x10x0x1 : tail0=1'b0;
        16'b0x0x11110x10x0x1 : tail0=1'b0;
        16'b110x11110x10x0x1 : tail0=1'b0;
        16'b10x111110x10x0x1 : tail0=1'b0;
        16'b0x1111110x10x0x1 : tail0=1'b0;
        16'b111111110x10x0x1 : tail0=1'b0;
        16'b10x0x0x0x110x0x1 : tail0=1'b0;
        16'b0x10x0x0x110x0x1 : tail0=1'b0;
        16'b1110x0x0x110x0x1 : tail0=1'b0;
        16'b0x0x10x0x110x0x1 : tail0=1'b0;
        16'b110x10x0x110x0x1 : tail0=1'b0;
        16'b10x110x0x110x0x1 : tail0=1'b0;
        16'b0x1110x0x110x0x1 : tail0=1'b0;
        16'b111110x0x110x0x1 : tail0=1'b0;
        16'b0x0x0x10x110x0x1 : tail0=1'b0;
        16'b110x0x10x110x0x1 : tail0=1'b0;
        16'b10x10x10x110x0x1 : tail0=1'b0;
        16'b0x110x10x110x0x1 : tail0=1'b0;
        16'b11110x10x110x0x1 : tail0=1'b0;
        16'b10x0x110x110x0x1 : tail0=1'b0;
        16'b0x10x110x110x0x1 : tail0=1'b0;
        16'b1110x110x110x0x1 : tail0=1'b0;
        16'b0x0x1110x110x0x1 : tail0=1'b0;
        16'b110x1110x110x0x1 : tail0=1'b0;
        16'b10x11110x110x0x1 : tail0=1'b0;
        16'b0x111110x110x0x1 : tail0=1'b0;
        16'b11111110x110x0x1 : tail0=1'b0;
        16'b0x0x0x0x1110x0x1 : tail0=1'b0;
        16'b110x0x0x1110x0x1 : tail0=1'b0;
        16'b10x10x0x1110x0x1 : tail0=1'b0;
        16'b0x110x0x1110x0x1 : tail0=1'b0;
        16'b11110x0x1110x0x1 : tail0=1'b0;
        16'b10x0x10x1110x0x1 : tail0=1'b0;
        16'b0x10x10x1110x0x1 : tail0=1'b0;
        16'b1110x10x1110x0x1 : tail0=1'b0;
        16'b0x0x110x1110x0x1 : tail0=1'b0;
        16'b110x110x1110x0x1 : tail0=1'b0;
        16'b10x1110x1110x0x1 : tail0=1'b0;
        16'b0x11110x1110x0x1 : tail0=1'b0;
        16'b1111110x1110x0x1 : tail0=1'b0;
        16'b10x0x0x11110x0x1 : tail0=1'b0;
        16'b0x10x0x11110x0x1 : tail0=1'b0;
        16'b1110x0x11110x0x1 : tail0=1'b0;
        16'b0x0x10x11110x0x1 : tail0=1'b0;
        16'b110x10x11110x0x1 : tail0=1'b0;
        16'b10x110x11110x0x1 : tail0=1'b0;
        16'b0x1110x11110x0x1 : tail0=1'b0;
        16'b111110x11110x0x1 : tail0=1'b0;
        16'b0x0x0x111110x0x1 : tail0=1'b0;
        16'b110x0x111110x0x1 : tail0=1'b0;
        16'b10x10x111110x0x1 : tail0=1'b0;
        16'b0x110x111110x0x1 : tail0=1'b0;
        16'b11110x111110x0x1 : tail0=1'b0;
        16'b10x0x1111110x0x1 : tail0=1'b0;
        16'b0x10x1111110x0x1 : tail0=1'b0;
        16'b1110x1111110x0x1 : tail0=1'b0;
        16'b0x0x11111110x0x1 : tail0=1'b0;
        16'b110x11111110x0x1 : tail0=1'b0;
        16'b10x111111110x0x1 : tail0=1'b0;
        16'b0x1111111110x0x1 : tail0=1'b0;
        16'b111111111110x0x1 : tail0=1'b0;
        16'b0x0x0x0x0x0x10x1 : tail0=1'b0;
        16'b110x0x0x0x0x10x1 : tail0=1'b0;
        16'b10x10x0x0x0x10x1 : tail0=1'b0;
        16'b0x110x0x0x0x10x1 : tail0=1'b0;
        16'b11110x0x0x0x10x1 : tail0=1'b0;
        16'b10x0x10x0x0x10x1 : tail0=1'b0;
        16'b0x10x10x0x0x10x1 : tail0=1'b0;
        16'b1110x10x0x0x10x1 : tail0=1'b0;
        16'b0x0x110x0x0x10x1 : tail0=1'b0;
        16'b110x110x0x0x10x1 : tail0=1'b0;
        16'b10x1110x0x0x10x1 : tail0=1'b0;
        16'b0x11110x0x0x10x1 : tail0=1'b0;
        16'b1111110x0x0x10x1 : tail0=1'b0;
        16'b10x0x0x10x0x10x1 : tail0=1'b0;
        16'b0x10x0x10x0x10x1 : tail0=1'b0;
        16'b1110x0x10x0x10x1 : tail0=1'b0;
        16'b0x0x10x10x0x10x1 : tail0=1'b0;
        16'b110x10x10x0x10x1 : tail0=1'b0;
        16'b10x110x10x0x10x1 : tail0=1'b0;
        16'b0x1110x10x0x10x1 : tail0=1'b0;
        16'b111110x10x0x10x1 : tail0=1'b0;
        16'b0x0x0x110x0x10x1 : tail0=1'b0;
        16'b110x0x110x0x10x1 : tail0=1'b0;
        16'b10x10x110x0x10x1 : tail0=1'b0;
        16'b0x110x110x0x10x1 : tail0=1'b0;
        16'b11110x110x0x10x1 : tail0=1'b0;
        16'b10x0x1110x0x10x1 : tail0=1'b0;
        16'b0x10x1110x0x10x1 : tail0=1'b0;
        16'b1110x1110x0x10x1 : tail0=1'b0;
        16'b0x0x11110x0x10x1 : tail0=1'b0;
        16'b110x11110x0x10x1 : tail0=1'b0;
        16'b10x111110x0x10x1 : tail0=1'b0;
        16'b0x1111110x0x10x1 : tail0=1'b0;
        16'b111111110x0x10x1 : tail0=1'b0;
        16'b10x0x0x0x10x10x1 : tail0=1'b0;
        16'b0x10x0x0x10x10x1 : tail0=1'b0;
        16'b1110x0x0x10x10x1 : tail0=1'b0;
        16'b0x0x10x0x10x10x1 : tail0=1'b0;
        16'b110x10x0x10x10x1 : tail0=1'b0;
        16'b10x110x0x10x10x1 : tail0=1'b0;
        16'b0x1110x0x10x10x1 : tail0=1'b0;
        16'b111110x0x10x10x1 : tail0=1'b0;
        16'b0x0x0x10x10x10x1 : tail0=1'b0;
        16'b110x0x10x10x10x1 : tail0=1'b0;
        16'b10x10x10x10x10x1 : tail0=1'b0;
        16'b0x110x10x10x10x1 : tail0=1'b0;
        16'b11110x10x10x10x1 : tail0=1'b0;
        16'b10x0x110x10x10x1 : tail0=1'b0;
        16'b0x10x110x10x10x1 : tail0=1'b0;
        16'b1110x110x10x10x1 : tail0=1'b0;
        16'b0x0x1110x10x10x1 : tail0=1'b0;
        16'b110x1110x10x10x1 : tail0=1'b0;
        16'b10x11110x10x10x1 : tail0=1'b0;
        16'b0x111110x10x10x1 : tail0=1'b0;
        16'b11111110x10x10x1 : tail0=1'b0;
        16'b0x0x0x0x110x10x1 : tail0=1'b0;
        16'b110x0x0x110x10x1 : tail0=1'b0;
        16'b10x10x0x110x10x1 : tail0=1'b0;
        16'b0x110x0x110x10x1 : tail0=1'b0;
        16'b11110x0x110x10x1 : tail0=1'b0;
        16'b10x0x10x110x10x1 : tail0=1'b0;
        16'b0x10x10x110x10x1 : tail0=1'b0;
        16'b1110x10x110x10x1 : tail0=1'b0;
        16'b0x0x110x110x10x1 : tail0=1'b0;
        16'b110x110x110x10x1 : tail0=1'b0;
        16'b10x1110x110x10x1 : tail0=1'b0;
        16'b0x11110x110x10x1 : tail0=1'b0;
        16'b1111110x110x10x1 : tail0=1'b0;
        16'b10x0x0x1110x10x1 : tail0=1'b0;
        16'b0x10x0x1110x10x1 : tail0=1'b0;
        16'b1110x0x1110x10x1 : tail0=1'b0;
        16'b0x0x10x1110x10x1 : tail0=1'b0;
        16'b110x10x1110x10x1 : tail0=1'b0;
        16'b10x110x1110x10x1 : tail0=1'b0;
        16'b0x1110x1110x10x1 : tail0=1'b0;
        16'b111110x1110x10x1 : tail0=1'b0;
        16'b0x0x0x11110x10x1 : tail0=1'b0;
        16'b110x0x11110x10x1 : tail0=1'b0;
        16'b10x10x11110x10x1 : tail0=1'b0;
        16'b0x110x11110x10x1 : tail0=1'b0;
        16'b11110x11110x10x1 : tail0=1'b0;
        16'b10x0x111110x10x1 : tail0=1'b0;
        16'b0x10x111110x10x1 : tail0=1'b0;
        16'b1110x111110x10x1 : tail0=1'b0;
        16'b0x0x1111110x10x1 : tail0=1'b0;
        16'b110x1111110x10x1 : tail0=1'b0;
        16'b10x11111110x10x1 : tail0=1'b0;
        16'b0x111111110x10x1 : tail0=1'b0;
        16'b11111111110x10x1 : tail0=1'b0;
        16'b10x0x0x0x0x110x1 : tail0=1'b0;
        16'b0x10x0x0x0x110x1 : tail0=1'b0;
        16'b1110x0x0x0x110x1 : tail0=1'b0;
        16'b0x0x10x0x0x110x1 : tail0=1'b0;
        16'b110x10x0x0x110x1 : tail0=1'b0;
        16'b10x110x0x0x110x1 : tail0=1'b0;
        16'b0x1110x0x0x110x1 : tail0=1'b0;
        16'b111110x0x0x110x1 : tail0=1'b0;
        16'b0x0x0x10x0x110x1 : tail0=1'b0;
        16'b110x0x10x0x110x1 : tail0=1'b0;
        16'b10x10x10x0x110x1 : tail0=1'b0;
        16'b0x110x10x0x110x1 : tail0=1'b0;
        16'b11110x10x0x110x1 : tail0=1'b0;
        16'b10x0x110x0x110x1 : tail0=1'b0;
        16'b0x10x110x0x110x1 : tail0=1'b0;
        16'b1110x110x0x110x1 : tail0=1'b0;
        16'b0x0x1110x0x110x1 : tail0=1'b0;
        16'b110x1110x0x110x1 : tail0=1'b0;
        16'b10x11110x0x110x1 : tail0=1'b0;
        16'b0x111110x0x110x1 : tail0=1'b0;
        16'b11111110x0x110x1 : tail0=1'b0;
        16'b0x0x0x0x10x110x1 : tail0=1'b0;
        16'b110x0x0x10x110x1 : tail0=1'b0;
        16'b10x10x0x10x110x1 : tail0=1'b0;
        16'b0x110x0x10x110x1 : tail0=1'b0;
        16'b11110x0x10x110x1 : tail0=1'b0;
        16'b10x0x10x10x110x1 : tail0=1'b0;
        16'b0x10x10x10x110x1 : tail0=1'b0;
        16'b1110x10x10x110x1 : tail0=1'b0;
        16'b0x0x110x10x110x1 : tail0=1'b0;
        16'b110x110x10x110x1 : tail0=1'b0;
        16'b10x1110x10x110x1 : tail0=1'b0;
        16'b0x11110x10x110x1 : tail0=1'b0;
        16'b1111110x10x110x1 : tail0=1'b0;
        16'b10x0x0x110x110x1 : tail0=1'b0;
        16'b0x10x0x110x110x1 : tail0=1'b0;
        16'b1110x0x110x110x1 : tail0=1'b0;
        16'b0x0x10x110x110x1 : tail0=1'b0;
        16'b110x10x110x110x1 : tail0=1'b0;
        16'b10x110x110x110x1 : tail0=1'b0;
        16'b0x1110x110x110x1 : tail0=1'b0;
        16'b111110x110x110x1 : tail0=1'b0;
        16'b0x0x0x1110x110x1 : tail0=1'b0;
        16'b110x0x1110x110x1 : tail0=1'b0;
        16'b10x10x1110x110x1 : tail0=1'b0;
        16'b0x110x1110x110x1 : tail0=1'b0;
        16'b11110x1110x110x1 : tail0=1'b0;
        16'b10x0x11110x110x1 : tail0=1'b0;
        16'b0x10x11110x110x1 : tail0=1'b0;
        16'b1110x11110x110x1 : tail0=1'b0;
        16'b0x0x111110x110x1 : tail0=1'b0;
        16'b110x111110x110x1 : tail0=1'b0;
        16'b10x1111110x110x1 : tail0=1'b0;
        16'b0x11111110x110x1 : tail0=1'b0;
        16'b1111111110x110x1 : tail0=1'b0;
        16'b0x0x0x0x0x1110x1 : tail0=1'b0;
        16'b110x0x0x0x1110x1 : tail0=1'b0;
        16'b10x10x0x0x1110x1 : tail0=1'b0;
        16'b0x110x0x0x1110x1 : tail0=1'b0;
        16'b11110x0x0x1110x1 : tail0=1'b0;
        16'b10x0x10x0x1110x1 : tail0=1'b0;
        16'b0x10x10x0x1110x1 : tail0=1'b0;
        16'b1110x10x0x1110x1 : tail0=1'b0;
        16'b0x0x110x0x1110x1 : tail0=1'b0;
        16'b110x110x0x1110x1 : tail0=1'b0;
        16'b10x1110x0x1110x1 : tail0=1'b0;
        16'b0x11110x0x1110x1 : tail0=1'b0;
        16'b1111110x0x1110x1 : tail0=1'b0;
        16'b10x0x0x10x1110x1 : tail0=1'b0;
        16'b0x10x0x10x1110x1 : tail0=1'b0;
        16'b1110x0x10x1110x1 : tail0=1'b0;
        16'b0x0x10x10x1110x1 : tail0=1'b0;
        16'b110x10x10x1110x1 : tail0=1'b0;
        16'b10x110x10x1110x1 : tail0=1'b0;
        16'b0x1110x10x1110x1 : tail0=1'b0;
        16'b111110x10x1110x1 : tail0=1'b0;
        16'b0x0x0x110x1110x1 : tail0=1'b0;
        16'b110x0x110x1110x1 : tail0=1'b0;
        16'b10x10x110x1110x1 : tail0=1'b0;
        16'b0x110x110x1110x1 : tail0=1'b0;
        16'b11110x110x1110x1 : tail0=1'b0;
        16'b10x0x1110x1110x1 : tail0=1'b0;
        16'b0x10x1110x1110x1 : tail0=1'b0;
        16'b1110x1110x1110x1 : tail0=1'b0;
        16'b0x0x11110x1110x1 : tail0=1'b0;
        16'b110x11110x1110x1 : tail0=1'b0;
        16'b10x111110x1110x1 : tail0=1'b0;
        16'b0x1111110x1110x1 : tail0=1'b0;
        16'b111111110x1110x1 : tail0=1'b0;
        16'b10x0x0x0x11110x1 : tail0=1'b0;
        16'b0x10x0x0x11110x1 : tail0=1'b0;
        16'b1110x0x0x11110x1 : tail0=1'b0;
        16'b0x0x10x0x11110x1 : tail0=1'b0;
        16'b110x10x0x11110x1 : tail0=1'b0;
        16'b10x110x0x11110x1 : tail0=1'b0;
        16'b0x1110x0x11110x1 : tail0=1'b0;
        16'b111110x0x11110x1 : tail0=1'b0;
        16'b0x0x0x10x11110x1 : tail0=1'b0;
        16'b110x0x10x11110x1 : tail0=1'b0;
        16'b10x10x10x11110x1 : tail0=1'b0;
        16'b0x110x10x11110x1 : tail0=1'b0;
        16'b11110x10x11110x1 : tail0=1'b0;
        16'b10x0x110x11110x1 : tail0=1'b0;
        16'b0x10x110x11110x1 : tail0=1'b0;
        16'b1110x110x11110x1 : tail0=1'b0;
        16'b0x0x1110x11110x1 : tail0=1'b0;
        16'b110x1110x11110x1 : tail0=1'b0;
        16'b10x11110x11110x1 : tail0=1'b0;
        16'b0x111110x11110x1 : tail0=1'b0;
        16'b11111110x11110x1 : tail0=1'b0;
        16'b0x0x0x0x111110x1 : tail0=1'b0;
        16'b110x0x0x111110x1 : tail0=1'b0;
        16'b10x10x0x111110x1 : tail0=1'b0;
        16'b0x110x0x111110x1 : tail0=1'b0;
        16'b11110x0x111110x1 : tail0=1'b0;
        16'b10x0x10x111110x1 : tail0=1'b0;
        16'b0x10x10x111110x1 : tail0=1'b0;
        16'b1110x10x111110x1 : tail0=1'b0;
        16'b0x0x110x111110x1 : tail0=1'b0;
        16'b110x110x111110x1 : tail0=1'b0;
        16'b10x1110x111110x1 : tail0=1'b0;
        16'b0x11110x111110x1 : tail0=1'b0;
        16'b1111110x111110x1 : tail0=1'b0;
        16'b10x0x0x1111110x1 : tail0=1'b0;
        16'b0x10x0x1111110x1 : tail0=1'b0;
        16'b1110x0x1111110x1 : tail0=1'b0;
        16'b0x0x10x1111110x1 : tail0=1'b0;
        16'b110x10x1111110x1 : tail0=1'b0;
        16'b10x110x1111110x1 : tail0=1'b0;
        16'b0x1110x1111110x1 : tail0=1'b0;
        16'b111110x1111110x1 : tail0=1'b0;
        16'b0x0x0x11111110x1 : tail0=1'b0;
        16'b110x0x11111110x1 : tail0=1'b0;
        16'b10x10x11111110x1 : tail0=1'b0;
        16'b0x110x11111110x1 : tail0=1'b0;
        16'b11110x11111110x1 : tail0=1'b0;
        16'b10x0x111111110x1 : tail0=1'b0;
        16'b0x10x111111110x1 : tail0=1'b0;
        16'b1110x111111110x1 : tail0=1'b0;
        16'b0x0x1111111110x1 : tail0=1'b0;
        16'b110x1111111110x1 : tail0=1'b0;
        16'b10x11111111110x1 : tail0=1'b0;
        16'b0x111111111110x1 : tail0=1'b0;
        16'b11111111111110x1 : tail0=1'b0;
        16'b0x0x0x0x0x0x0x11 : tail0=1'b0;
        16'b110x0x0x0x0x0x11 : tail0=1'b0;
        16'b10x10x0x0x0x0x11 : tail0=1'b0;
        16'b0x110x0x0x0x0x11 : tail0=1'b0;
        16'b11110x0x0x0x0x11 : tail0=1'b0;
        16'b10x0x10x0x0x0x11 : tail0=1'b0;
        16'b0x10x10x0x0x0x11 : tail0=1'b0;
        16'b1110x10x0x0x0x11 : tail0=1'b0;
        16'b0x0x110x0x0x0x11 : tail0=1'b0;
        16'b110x110x0x0x0x11 : tail0=1'b0;
        16'b10x1110x0x0x0x11 : tail0=1'b0;
        16'b0x11110x0x0x0x11 : tail0=1'b0;
        16'b1111110x0x0x0x11 : tail0=1'b0;
        16'b10x0x0x10x0x0x11 : tail0=1'b0;
        16'b0x10x0x10x0x0x11 : tail0=1'b0;
        16'b1110x0x10x0x0x11 : tail0=1'b0;
        16'b0x0x10x10x0x0x11 : tail0=1'b0;
        16'b110x10x10x0x0x11 : tail0=1'b0;
        16'b10x110x10x0x0x11 : tail0=1'b0;
        16'b0x1110x10x0x0x11 : tail0=1'b0;
        16'b111110x10x0x0x11 : tail0=1'b0;
        16'b0x0x0x110x0x0x11 : tail0=1'b0;
        16'b110x0x110x0x0x11 : tail0=1'b0;
        16'b10x10x110x0x0x11 : tail0=1'b0;
        16'b0x110x110x0x0x11 : tail0=1'b0;
        16'b11110x110x0x0x11 : tail0=1'b0;
        16'b10x0x1110x0x0x11 : tail0=1'b0;
        16'b0x10x1110x0x0x11 : tail0=1'b0;
        16'b1110x1110x0x0x11 : tail0=1'b0;
        16'b0x0x11110x0x0x11 : tail0=1'b0;
        16'b110x11110x0x0x11 : tail0=1'b0;
        16'b10x111110x0x0x11 : tail0=1'b0;
        16'b0x1111110x0x0x11 : tail0=1'b0;
        16'b111111110x0x0x11 : tail0=1'b0;
        16'b10x0x0x0x10x0x11 : tail0=1'b0;
        16'b0x10x0x0x10x0x11 : tail0=1'b0;
        16'b1110x0x0x10x0x11 : tail0=1'b0;
        16'b0x0x10x0x10x0x11 : tail0=1'b0;
        16'b110x10x0x10x0x11 : tail0=1'b0;
        16'b10x110x0x10x0x11 : tail0=1'b0;
        16'b0x1110x0x10x0x11 : tail0=1'b0;
        16'b111110x0x10x0x11 : tail0=1'b0;
        16'b0x0x0x10x10x0x11 : tail0=1'b0;
        16'b110x0x10x10x0x11 : tail0=1'b0;
        16'b10x10x10x10x0x11 : tail0=1'b0;
        16'b0x110x10x10x0x11 : tail0=1'b0;
        16'b11110x10x10x0x11 : tail0=1'b0;
        16'b10x0x110x10x0x11 : tail0=1'b0;
        16'b0x10x110x10x0x11 : tail0=1'b0;
        16'b1110x110x10x0x11 : tail0=1'b0;
        16'b0x0x1110x10x0x11 : tail0=1'b0;
        16'b110x1110x10x0x11 : tail0=1'b0;
        16'b10x11110x10x0x11 : tail0=1'b0;
        16'b0x111110x10x0x11 : tail0=1'b0;
        16'b11111110x10x0x11 : tail0=1'b0;
        16'b0x0x0x0x110x0x11 : tail0=1'b0;
        16'b110x0x0x110x0x11 : tail0=1'b0;
        16'b10x10x0x110x0x11 : tail0=1'b0;
        16'b0x110x0x110x0x11 : tail0=1'b0;
        16'b11110x0x110x0x11 : tail0=1'b0;
        16'b10x0x10x110x0x11 : tail0=1'b0;
        16'b0x10x10x110x0x11 : tail0=1'b0;
        16'b1110x10x110x0x11 : tail0=1'b0;
        16'b0x0x110x110x0x11 : tail0=1'b0;
        16'b110x110x110x0x11 : tail0=1'b0;
        16'b10x1110x110x0x11 : tail0=1'b0;
        16'b0x11110x110x0x11 : tail0=1'b0;
        16'b1111110x110x0x11 : tail0=1'b0;
        16'b10x0x0x1110x0x11 : tail0=1'b0;
        16'b0x10x0x1110x0x11 : tail0=1'b0;
        16'b1110x0x1110x0x11 : tail0=1'b0;
        16'b0x0x10x1110x0x11 : tail0=1'b0;
        16'b110x10x1110x0x11 : tail0=1'b0;
        16'b10x110x1110x0x11 : tail0=1'b0;
        16'b0x1110x1110x0x11 : tail0=1'b0;
        16'b111110x1110x0x11 : tail0=1'b0;
        16'b0x0x0x11110x0x11 : tail0=1'b0;
        16'b110x0x11110x0x11 : tail0=1'b0;
        16'b10x10x11110x0x11 : tail0=1'b0;
        16'b0x110x11110x0x11 : tail0=1'b0;
        16'b11110x11110x0x11 : tail0=1'b0;
        16'b10x0x111110x0x11 : tail0=1'b0;
        16'b0x10x111110x0x11 : tail0=1'b0;
        16'b1110x111110x0x11 : tail0=1'b0;
        16'b0x0x1111110x0x11 : tail0=1'b0;
        16'b110x1111110x0x11 : tail0=1'b0;
        16'b10x11111110x0x11 : tail0=1'b0;
        16'b0x111111110x0x11 : tail0=1'b0;
        16'b11111111110x0x11 : tail0=1'b0;
        16'b10x0x0x0x0x10x11 : tail0=1'b0;
        16'b0x10x0x0x0x10x11 : tail0=1'b0;
        16'b1110x0x0x0x10x11 : tail0=1'b0;
        16'b0x0x10x0x0x10x11 : tail0=1'b0;
        16'b110x10x0x0x10x11 : tail0=1'b0;
        16'b10x110x0x0x10x11 : tail0=1'b0;
        16'b0x1110x0x0x10x11 : tail0=1'b0;
        16'b111110x0x0x10x11 : tail0=1'b0;
        16'b0x0x0x10x0x10x11 : tail0=1'b0;
        16'b110x0x10x0x10x11 : tail0=1'b0;
        16'b10x10x10x0x10x11 : tail0=1'b0;
        16'b0x110x10x0x10x11 : tail0=1'b0;
        16'b11110x10x0x10x11 : tail0=1'b0;
        16'b10x0x110x0x10x11 : tail0=1'b0;
        16'b0x10x110x0x10x11 : tail0=1'b0;
        16'b1110x110x0x10x11 : tail0=1'b0;
        16'b0x0x1110x0x10x11 : tail0=1'b0;
        16'b110x1110x0x10x11 : tail0=1'b0;
        16'b10x11110x0x10x11 : tail0=1'b0;
        16'b0x111110x0x10x11 : tail0=1'b0;
        16'b11111110x0x10x11 : tail0=1'b0;
        16'b0x0x0x0x10x10x11 : tail0=1'b0;
        16'b110x0x0x10x10x11 : tail0=1'b0;
        16'b10x10x0x10x10x11 : tail0=1'b0;
        16'b0x110x0x10x10x11 : tail0=1'b0;
        16'b11110x0x10x10x11 : tail0=1'b0;
        16'b10x0x10x10x10x11 : tail0=1'b0;
        16'b0x10x10x10x10x11 : tail0=1'b0;
        16'b1110x10x10x10x11 : tail0=1'b0;
        16'b0x0x110x10x10x11 : tail0=1'b0;
        16'b110x110x10x10x11 : tail0=1'b0;
        16'b10x1110x10x10x11 : tail0=1'b0;
        16'b0x11110x10x10x11 : tail0=1'b0;
        16'b1111110x10x10x11 : tail0=1'b0;
        16'b10x0x0x110x10x11 : tail0=1'b0;
        16'b0x10x0x110x10x11 : tail0=1'b0;
        16'b1110x0x110x10x11 : tail0=1'b0;
        16'b0x0x10x110x10x11 : tail0=1'b0;
        16'b110x10x110x10x11 : tail0=1'b0;
        16'b10x110x110x10x11 : tail0=1'b0;
        16'b0x1110x110x10x11 : tail0=1'b0;
        16'b111110x110x10x11 : tail0=1'b0;
        16'b0x0x0x1110x10x11 : tail0=1'b0;
        16'b110x0x1110x10x11 : tail0=1'b0;
        16'b10x10x1110x10x11 : tail0=1'b0;
        16'b0x110x1110x10x11 : tail0=1'b0;
        16'b11110x1110x10x11 : tail0=1'b0;
        16'b10x0x11110x10x11 : tail0=1'b0;
        16'b0x10x11110x10x11 : tail0=1'b0;
        16'b1110x11110x10x11 : tail0=1'b0;
        16'b0x0x111110x10x11 : tail0=1'b0;
        16'b110x111110x10x11 : tail0=1'b0;
        16'b10x1111110x10x11 : tail0=1'b0;
        16'b0x11111110x10x11 : tail0=1'b0;
        16'b1111111110x10x11 : tail0=1'b0;
        16'b0x0x0x0x0x110x11 : tail0=1'b0;
        16'b110x0x0x0x110x11 : tail0=1'b0;
        16'b10x10x0x0x110x11 : tail0=1'b0;
        16'b0x110x0x0x110x11 : tail0=1'b0;
        16'b11110x0x0x110x11 : tail0=1'b0;
        16'b10x0x10x0x110x11 : tail0=1'b0;
        16'b0x10x10x0x110x11 : tail0=1'b0;
        16'b1110x10x0x110x11 : tail0=1'b0;
        16'b0x0x110x0x110x11 : tail0=1'b0;
        16'b110x110x0x110x11 : tail0=1'b0;
        16'b10x1110x0x110x11 : tail0=1'b0;
        16'b0x11110x0x110x11 : tail0=1'b0;
        16'b1111110x0x110x11 : tail0=1'b0;
        16'b10x0x0x10x110x11 : tail0=1'b0;
        16'b0x10x0x10x110x11 : tail0=1'b0;
        16'b1110x0x10x110x11 : tail0=1'b0;
        16'b0x0x10x10x110x11 : tail0=1'b0;
        16'b110x10x10x110x11 : tail0=1'b0;
        16'b10x110x10x110x11 : tail0=1'b0;
        16'b0x1110x10x110x11 : tail0=1'b0;
        16'b111110x10x110x11 : tail0=1'b0;
        16'b0x0x0x110x110x11 : tail0=1'b0;
        16'b110x0x110x110x11 : tail0=1'b0;
        16'b10x10x110x110x11 : tail0=1'b0;
        16'b0x110x110x110x11 : tail0=1'b0;
        16'b11110x110x110x11 : tail0=1'b0;
        16'b10x0x1110x110x11 : tail0=1'b0;
        16'b0x10x1110x110x11 : tail0=1'b0;
        16'b1110x1110x110x11 : tail0=1'b0;
        16'b0x0x11110x110x11 : tail0=1'b0;
        16'b110x11110x110x11 : tail0=1'b0;
        16'b10x111110x110x11 : tail0=1'b0;
        16'b0x1111110x110x11 : tail0=1'b0;
        16'b111111110x110x11 : tail0=1'b0;
        16'b10x0x0x0x1110x11 : tail0=1'b0;
        16'b0x10x0x0x1110x11 : tail0=1'b0;
        16'b1110x0x0x1110x11 : tail0=1'b0;
        16'b0x0x10x0x1110x11 : tail0=1'b0;
        16'b110x10x0x1110x11 : tail0=1'b0;
        16'b10x110x0x1110x11 : tail0=1'b0;
        16'b0x1110x0x1110x11 : tail0=1'b0;
        16'b111110x0x1110x11 : tail0=1'b0;
        16'b0x0x0x10x1110x11 : tail0=1'b0;
        16'b110x0x10x1110x11 : tail0=1'b0;
        16'b10x10x10x1110x11 : tail0=1'b0;
        16'b0x110x10x1110x11 : tail0=1'b0;
        16'b11110x10x1110x11 : tail0=1'b0;
        16'b10x0x110x1110x11 : tail0=1'b0;
        16'b0x10x110x1110x11 : tail0=1'b0;
        16'b1110x110x1110x11 : tail0=1'b0;
        16'b0x0x1110x1110x11 : tail0=1'b0;
        16'b110x1110x1110x11 : tail0=1'b0;
        16'b10x11110x1110x11 : tail0=1'b0;
        16'b0x111110x1110x11 : tail0=1'b0;
        16'b11111110x1110x11 : tail0=1'b0;
        16'b0x0x0x0x11110x11 : tail0=1'b0;
        16'b110x0x0x11110x11 : tail0=1'b0;
        16'b10x10x0x11110x11 : tail0=1'b0;
        16'b0x110x0x11110x11 : tail0=1'b0;
        16'b11110x0x11110x11 : tail0=1'b0;
        16'b10x0x10x11110x11 : tail0=1'b0;
        16'b0x10x10x11110x11 : tail0=1'b0;
        16'b1110x10x11110x11 : tail0=1'b0;
        16'b0x0x110x11110x11 : tail0=1'b0;
        16'b110x110x11110x11 : tail0=1'b0;
        16'b10x1110x11110x11 : tail0=1'b0;
        16'b0x11110x11110x11 : tail0=1'b0;
        16'b1111110x11110x11 : tail0=1'b0;
        16'b10x0x0x111110x11 : tail0=1'b0;
        16'b0x10x0x111110x11 : tail0=1'b0;
        16'b1110x0x111110x11 : tail0=1'b0;
        16'b0x0x10x111110x11 : tail0=1'b0;
        16'b110x10x111110x11 : tail0=1'b0;
        16'b10x110x111110x11 : tail0=1'b0;
        16'b0x1110x111110x11 : tail0=1'b0;
        16'b111110x111110x11 : tail0=1'b0;
        16'b0x0x0x1111110x11 : tail0=1'b0;
        16'b110x0x1111110x11 : tail0=1'b0;
        16'b10x10x1111110x11 : tail0=1'b0;
        16'b0x110x1111110x11 : tail0=1'b0;
        16'b11110x1111110x11 : tail0=1'b0;
        16'b10x0x11111110x11 : tail0=1'b0;
        16'b0x10x11111110x11 : tail0=1'b0;
        16'b1110x11111110x11 : tail0=1'b0;
        16'b0x0x111111110x11 : tail0=1'b0;
        16'b110x111111110x11 : tail0=1'b0;
        16'b10x1111111110x11 : tail0=1'b0;
        16'b0x11111111110x11 : tail0=1'b0;
        16'b1111111111110x11 : tail0=1'b0;
        16'b10x0x0x0x0x0x111 : tail0=1'b0;
        16'b0x10x0x0x0x0x111 : tail0=1'b0;
        16'b1110x0x0x0x0x111 : tail0=1'b0;
        16'b0x0x10x0x0x0x111 : tail0=1'b0;
        16'b110x10x0x0x0x111 : tail0=1'b0;
        16'b10x110x0x0x0x111 : tail0=1'b0;
        16'b0x1110x0x0x0x111 : tail0=1'b0;
        16'b111110x0x0x0x111 : tail0=1'b0;
        16'b0x0x0x10x0x0x111 : tail0=1'b0;
        16'b110x0x10x0x0x111 : tail0=1'b0;
        16'b10x10x10x0x0x111 : tail0=1'b0;
        16'b0x110x10x0x0x111 : tail0=1'b0;
        16'b11110x10x0x0x111 : tail0=1'b0;
        16'b10x0x110x0x0x111 : tail0=1'b0;
        16'b0x10x110x0x0x111 : tail0=1'b0;
        16'b1110x110x0x0x111 : tail0=1'b0;
        16'b0x0x1110x0x0x111 : tail0=1'b0;
        16'b110x1110x0x0x111 : tail0=1'b0;
        16'b10x11110x0x0x111 : tail0=1'b0;
        16'b0x111110x0x0x111 : tail0=1'b0;
        16'b11111110x0x0x111 : tail0=1'b0;
        16'b0x0x0x0x10x0x111 : tail0=1'b0;
        16'b110x0x0x10x0x111 : tail0=1'b0;
        16'b10x10x0x10x0x111 : tail0=1'b0;
        16'b0x110x0x10x0x111 : tail0=1'b0;
        16'b11110x0x10x0x111 : tail0=1'b0;
        16'b10x0x10x10x0x111 : tail0=1'b0;
        16'b0x10x10x10x0x111 : tail0=1'b0;
        16'b1110x10x10x0x111 : tail0=1'b0;
        16'b0x0x110x10x0x111 : tail0=1'b0;
        16'b110x110x10x0x111 : tail0=1'b0;
        16'b10x1110x10x0x111 : tail0=1'b0;
        16'b0x11110x10x0x111 : tail0=1'b0;
        16'b1111110x10x0x111 : tail0=1'b0;
        16'b10x0x0x110x0x111 : tail0=1'b0;
        16'b0x10x0x110x0x111 : tail0=1'b0;
        16'b1110x0x110x0x111 : tail0=1'b0;
        16'b0x0x10x110x0x111 : tail0=1'b0;
        16'b110x10x110x0x111 : tail0=1'b0;
        16'b10x110x110x0x111 : tail0=1'b0;
        16'b0x1110x110x0x111 : tail0=1'b0;
        16'b111110x110x0x111 : tail0=1'b0;
        16'b0x0x0x1110x0x111 : tail0=1'b0;
        16'b110x0x1110x0x111 : tail0=1'b0;
        16'b10x10x1110x0x111 : tail0=1'b0;
        16'b0x110x1110x0x111 : tail0=1'b0;
        16'b11110x1110x0x111 : tail0=1'b0;
        16'b10x0x11110x0x111 : tail0=1'b0;
        16'b0x10x11110x0x111 : tail0=1'b0;
        16'b1110x11110x0x111 : tail0=1'b0;
        16'b0x0x111110x0x111 : tail0=1'b0;
        16'b110x111110x0x111 : tail0=1'b0;
        16'b10x1111110x0x111 : tail0=1'b0;
        16'b0x11111110x0x111 : tail0=1'b0;
        16'b1111111110x0x111 : tail0=1'b0;
        16'b0x0x0x0x0x10x111 : tail0=1'b0;
        16'b110x0x0x0x10x111 : tail0=1'b0;
        16'b10x10x0x0x10x111 : tail0=1'b0;
        16'b0x110x0x0x10x111 : tail0=1'b0;
        16'b11110x0x0x10x111 : tail0=1'b0;
        16'b10x0x10x0x10x111 : tail0=1'b0;
        16'b0x10x10x0x10x111 : tail0=1'b0;
        16'b1110x10x0x10x111 : tail0=1'b0;
        16'b0x0x110x0x10x111 : tail0=1'b0;
        16'b110x110x0x10x111 : tail0=1'b0;
        16'b10x1110x0x10x111 : tail0=1'b0;
        16'b0x11110x0x10x111 : tail0=1'b0;
        16'b1111110x0x10x111 : tail0=1'b0;
        16'b10x0x0x10x10x111 : tail0=1'b0;
        16'b0x10x0x10x10x111 : tail0=1'b0;
        16'b1110x0x10x10x111 : tail0=1'b0;
        16'b0x0x10x10x10x111 : tail0=1'b0;
        16'b110x10x10x10x111 : tail0=1'b0;
        16'b10x110x10x10x111 : tail0=1'b0;
        16'b0x1110x10x10x111 : tail0=1'b0;
        16'b111110x10x10x111 : tail0=1'b0;
        16'b0x0x0x110x10x111 : tail0=1'b0;
        16'b110x0x110x10x111 : tail0=1'b0;
        16'b10x10x110x10x111 : tail0=1'b0;
        16'b0x110x110x10x111 : tail0=1'b0;
        16'b11110x110x10x111 : tail0=1'b0;
        16'b10x0x1110x10x111 : tail0=1'b0;
        16'b0x10x1110x10x111 : tail0=1'b0;
        16'b1110x1110x10x111 : tail0=1'b0;
        16'b0x0x11110x10x111 : tail0=1'b0;
        16'b110x11110x10x111 : tail0=1'b0;
        16'b10x111110x10x111 : tail0=1'b0;
        16'b0x1111110x10x111 : tail0=1'b0;
        16'b111111110x10x111 : tail0=1'b0;
        16'b10x0x0x0x110x111 : tail0=1'b0;
        16'b0x10x0x0x110x111 : tail0=1'b0;
        16'b1110x0x0x110x111 : tail0=1'b0;
        16'b0x0x10x0x110x111 : tail0=1'b0;
        16'b110x10x0x110x111 : tail0=1'b0;
        16'b10x110x0x110x111 : tail0=1'b0;
        16'b0x1110x0x110x111 : tail0=1'b0;
        16'b111110x0x110x111 : tail0=1'b0;
        16'b0x0x0x10x110x111 : tail0=1'b0;
        16'b110x0x10x110x111 : tail0=1'b0;
        16'b10x10x10x110x111 : tail0=1'b0;
        16'b0x110x10x110x111 : tail0=1'b0;
        16'b11110x10x110x111 : tail0=1'b0;
        16'b10x0x110x110x111 : tail0=1'b0;
        16'b0x10x110x110x111 : tail0=1'b0;
        16'b1110x110x110x111 : tail0=1'b0;
        16'b0x0x1110x110x111 : tail0=1'b0;
        16'b110x1110x110x111 : tail0=1'b0;
        16'b10x11110x110x111 : tail0=1'b0;
        16'b0x111110x110x111 : tail0=1'b0;
        16'b11111110x110x111 : tail0=1'b0;
        16'b0x0x0x0x1110x111 : tail0=1'b0;
        16'b110x0x0x1110x111 : tail0=1'b0;
        16'b10x10x0x1110x111 : tail0=1'b0;
        16'b0x110x0x1110x111 : tail0=1'b0;
        16'b11110x0x1110x111 : tail0=1'b0;
        16'b10x0x10x1110x111 : tail0=1'b0;
        16'b0x10x10x1110x111 : tail0=1'b0;
        16'b1110x10x1110x111 : tail0=1'b0;
        16'b0x0x110x1110x111 : tail0=1'b0;
        16'b110x110x1110x111 : tail0=1'b0;
        16'b10x1110x1110x111 : tail0=1'b0;
        16'b0x11110x1110x111 : tail0=1'b0;
        16'b1111110x1110x111 : tail0=1'b0;
        16'b10x0x0x11110x111 : tail0=1'b0;
        16'b0x10x0x11110x111 : tail0=1'b0;
        16'b1110x0x11110x111 : tail0=1'b0;
        16'b0x0x10x11110x111 : tail0=1'b0;
        16'b110x10x11110x111 : tail0=1'b0;
        16'b10x110x11110x111 : tail0=1'b0;
        16'b0x1110x11110x111 : tail0=1'b0;
        16'b111110x11110x111 : tail0=1'b0;
        16'b0x0x0x111110x111 : tail0=1'b0;
        16'b110x0x111110x111 : tail0=1'b0;
        16'b10x10x111110x111 : tail0=1'b0;
        16'b0x110x111110x111 : tail0=1'b0;
        16'b11110x111110x111 : tail0=1'b0;
        16'b10x0x1111110x111 : tail0=1'b0;
        16'b0x10x1111110x111 : tail0=1'b0;
        16'b1110x1111110x111 : tail0=1'b0;
        16'b0x0x11111110x111 : tail0=1'b0;
        16'b110x11111110x111 : tail0=1'b0;
        16'b10x111111110x111 : tail0=1'b0;
        16'b0x1111111110x111 : tail0=1'b0;
        16'b111111111110x111 : tail0=1'b0;
        16'b0x0x0x0x0x0x1111 : tail0=1'b0;
        16'b110x0x0x0x0x1111 : tail0=1'b0;
        16'b10x10x0x0x0x1111 : tail0=1'b0;
        16'b0x110x0x0x0x1111 : tail0=1'b0;
        16'b11110x0x0x0x1111 : tail0=1'b0;
        16'b10x0x10x0x0x1111 : tail0=1'b0;
        16'b0x10x10x0x0x1111 : tail0=1'b0;
        16'b1110x10x0x0x1111 : tail0=1'b0;
        16'b0x0x110x0x0x1111 : tail0=1'b0;
        16'b110x110x0x0x1111 : tail0=1'b0;
        16'b10x1110x0x0x1111 : tail0=1'b0;
        16'b0x11110x0x0x1111 : tail0=1'b0;
        16'b1111110x0x0x1111 : tail0=1'b0;
        16'b10x0x0x10x0x1111 : tail0=1'b0;
        16'b0x10x0x10x0x1111 : tail0=1'b0;
        16'b1110x0x10x0x1111 : tail0=1'b0;
        16'b0x0x10x10x0x1111 : tail0=1'b0;
        16'b110x10x10x0x1111 : tail0=1'b0;
        16'b10x110x10x0x1111 : tail0=1'b0;
        16'b0x1110x10x0x1111 : tail0=1'b0;
        16'b111110x10x0x1111 : tail0=1'b0;
        16'b0x0x0x110x0x1111 : tail0=1'b0;
        16'b110x0x110x0x1111 : tail0=1'b0;
        16'b10x10x110x0x1111 : tail0=1'b0;
        16'b0x110x110x0x1111 : tail0=1'b0;
        16'b11110x110x0x1111 : tail0=1'b0;
        16'b10x0x1110x0x1111 : tail0=1'b0;
        16'b0x10x1110x0x1111 : tail0=1'b0;
        16'b1110x1110x0x1111 : tail0=1'b0;
        16'b0x0x11110x0x1111 : tail0=1'b0;
        16'b110x11110x0x1111 : tail0=1'b0;
        16'b10x111110x0x1111 : tail0=1'b0;
        16'b0x1111110x0x1111 : tail0=1'b0;
        16'b111111110x0x1111 : tail0=1'b0;
        16'b10x0x0x0x10x1111 : tail0=1'b0;
        16'b0x10x0x0x10x1111 : tail0=1'b0;
        16'b1110x0x0x10x1111 : tail0=1'b0;
        16'b0x0x10x0x10x1111 : tail0=1'b0;
        16'b110x10x0x10x1111 : tail0=1'b0;
        16'b10x110x0x10x1111 : tail0=1'b0;
        16'b0x1110x0x10x1111 : tail0=1'b0;
        16'b111110x0x10x1111 : tail0=1'b0;
        16'b0x0x0x10x10x1111 : tail0=1'b0;
        16'b110x0x10x10x1111 : tail0=1'b0;
        16'b10x10x10x10x1111 : tail0=1'b0;
        16'b0x110x10x10x1111 : tail0=1'b0;
        16'b11110x10x10x1111 : tail0=1'b0;
        16'b10x0x110x10x1111 : tail0=1'b0;
        16'b0x10x110x10x1111 : tail0=1'b0;
        16'b1110x110x10x1111 : tail0=1'b0;
        16'b0x0x1110x10x1111 : tail0=1'b0;
        16'b110x1110x10x1111 : tail0=1'b0;
        16'b10x11110x10x1111 : tail0=1'b0;
        16'b0x111110x10x1111 : tail0=1'b0;
        16'b11111110x10x1111 : tail0=1'b0;
        16'b0x0x0x0x110x1111 : tail0=1'b0;
        16'b110x0x0x110x1111 : tail0=1'b0;
        16'b10x10x0x110x1111 : tail0=1'b0;
        16'b0x110x0x110x1111 : tail0=1'b0;
        16'b11110x0x110x1111 : tail0=1'b0;
        16'b10x0x10x110x1111 : tail0=1'b0;
        16'b0x10x10x110x1111 : tail0=1'b0;
        16'b1110x10x110x1111 : tail0=1'b0;
        16'b0x0x110x110x1111 : tail0=1'b0;
        16'b110x110x110x1111 : tail0=1'b0;
        16'b10x1110x110x1111 : tail0=1'b0;
        16'b0x11110x110x1111 : tail0=1'b0;
        16'b1111110x110x1111 : tail0=1'b0;
        16'b10x0x0x1110x1111 : tail0=1'b0;
        16'b0x10x0x1110x1111 : tail0=1'b0;
        16'b1110x0x1110x1111 : tail0=1'b0;
        16'b0x0x10x1110x1111 : tail0=1'b0;
        16'b110x10x1110x1111 : tail0=1'b0;
        16'b10x110x1110x1111 : tail0=1'b0;
        16'b0x1110x1110x1111 : tail0=1'b0;
        16'b111110x1110x1111 : tail0=1'b0;
        16'b0x0x0x11110x1111 : tail0=1'b0;
        16'b110x0x11110x1111 : tail0=1'b0;
        16'b10x10x11110x1111 : tail0=1'b0;
        16'b0x110x11110x1111 : tail0=1'b0;
        16'b11110x11110x1111 : tail0=1'b0;
        16'b10x0x111110x1111 : tail0=1'b0;
        16'b0x10x111110x1111 : tail0=1'b0;
        16'b1110x111110x1111 : tail0=1'b0;
        16'b0x0x1111110x1111 : tail0=1'b0;
        16'b110x1111110x1111 : tail0=1'b0;
        16'b10x11111110x1111 : tail0=1'b0;
        16'b0x111111110x1111 : tail0=1'b0;
        16'b11111111110x1111 : tail0=1'b0;
        16'b10x0x0x0x0x11111 : tail0=1'b0;
        16'b0x10x0x0x0x11111 : tail0=1'b0;
        16'b1110x0x0x0x11111 : tail0=1'b0;
        16'b0x0x10x0x0x11111 : tail0=1'b0;
        16'b110x10x0x0x11111 : tail0=1'b0;
        16'b10x110x0x0x11111 : tail0=1'b0;
        16'b0x1110x0x0x11111 : tail0=1'b0;
        16'b111110x0x0x11111 : tail0=1'b0;
        16'b0x0x0x10x0x11111 : tail0=1'b0;
        16'b110x0x10x0x11111 : tail0=1'b0;
        16'b10x10x10x0x11111 : tail0=1'b0;
        16'b0x110x10x0x11111 : tail0=1'b0;
        16'b11110x10x0x11111 : tail0=1'b0;
        16'b10x0x110x0x11111 : tail0=1'b0;
        16'b0x10x110x0x11111 : tail0=1'b0;
        16'b1110x110x0x11111 : tail0=1'b0;
        16'b0x0x1110x0x11111 : tail0=1'b0;
        16'b110x1110x0x11111 : tail0=1'b0;
        16'b10x11110x0x11111 : tail0=1'b0;
        16'b0x111110x0x11111 : tail0=1'b0;
        16'b11111110x0x11111 : tail0=1'b0;
        16'b0x0x0x0x10x11111 : tail0=1'b0;
        16'b110x0x0x10x11111 : tail0=1'b0;
        16'b10x10x0x10x11111 : tail0=1'b0;
        16'b0x110x0x10x11111 : tail0=1'b0;
        16'b11110x0x10x11111 : tail0=1'b0;
        16'b10x0x10x10x11111 : tail0=1'b0;
        16'b0x10x10x10x11111 : tail0=1'b0;
        16'b1110x10x10x11111 : tail0=1'b0;
        16'b0x0x110x10x11111 : tail0=1'b0;
        16'b110x110x10x11111 : tail0=1'b0;
        16'b10x1110x10x11111 : tail0=1'b0;
        16'b0x11110x10x11111 : tail0=1'b0;
        16'b1111110x10x11111 : tail0=1'b0;
        16'b10x0x0x110x11111 : tail0=1'b0;
        16'b0x10x0x110x11111 : tail0=1'b0;
        16'b1110x0x110x11111 : tail0=1'b0;
        16'b0x0x10x110x11111 : tail0=1'b0;
        16'b110x10x110x11111 : tail0=1'b0;
        16'b10x110x110x11111 : tail0=1'b0;
        16'b0x1110x110x11111 : tail0=1'b0;
        16'b111110x110x11111 : tail0=1'b0;
        16'b0x0x0x1110x11111 : tail0=1'b0;
        16'b110x0x1110x11111 : tail0=1'b0;
        16'b10x10x1110x11111 : tail0=1'b0;
        16'b0x110x1110x11111 : tail0=1'b0;
        16'b11110x1110x11111 : tail0=1'b0;
        16'b10x0x11110x11111 : tail0=1'b0;
        16'b0x10x11110x11111 : tail0=1'b0;
        16'b1110x11110x11111 : tail0=1'b0;
        16'b0x0x111110x11111 : tail0=1'b0;
        16'b110x111110x11111 : tail0=1'b0;
        16'b10x1111110x11111 : tail0=1'b0;
        16'b0x11111110x11111 : tail0=1'b0;
        16'b1111111110x11111 : tail0=1'b0;
        16'b0x0x0x0x0x111111 : tail0=1'b0;
        16'b110x0x0x0x111111 : tail0=1'b0;
        16'b10x10x0x0x111111 : tail0=1'b0;
        16'b0x110x0x0x111111 : tail0=1'b0;
        16'b11110x0x0x111111 : tail0=1'b0;
        16'b10x0x10x0x111111 : tail0=1'b0;
        16'b0x10x10x0x111111 : tail0=1'b0;
        16'b1110x10x0x111111 : tail0=1'b0;
        16'b0x0x110x0x111111 : tail0=1'b0;
        16'b110x110x0x111111 : tail0=1'b0;
        16'b10x1110x0x111111 : tail0=1'b0;
        16'b0x11110x0x111111 : tail0=1'b0;
        16'b1111110x0x111111 : tail0=1'b0;
        16'b10x0x0x10x111111 : tail0=1'b0;
        16'b0x10x0x10x111111 : tail0=1'b0;
        16'b1110x0x10x111111 : tail0=1'b0;
        16'b0x0x10x10x111111 : tail0=1'b0;
        16'b110x10x10x111111 : tail0=1'b0;
        16'b10x110x10x111111 : tail0=1'b0;
        16'b0x1110x10x111111 : tail0=1'b0;
        16'b111110x10x111111 : tail0=1'b0;
        16'b0x0x0x110x111111 : tail0=1'b0;
        16'b110x0x110x111111 : tail0=1'b0;
        16'b10x10x110x111111 : tail0=1'b0;
        16'b0x110x110x111111 : tail0=1'b0;
        16'b11110x110x111111 : tail0=1'b0;
        16'b10x0x1110x111111 : tail0=1'b0;
        16'b0x10x1110x111111 : tail0=1'b0;
        16'b1110x1110x111111 : tail0=1'b0;
        16'b0x0x11110x111111 : tail0=1'b0;
        16'b110x11110x111111 : tail0=1'b0;
        16'b10x111110x111111 : tail0=1'b0;
        16'b0x1111110x111111 : tail0=1'b0;
        16'b111111110x111111 : tail0=1'b0;
        16'b10x0x0x0x1111111 : tail0=1'b0;
        16'b0x10x0x0x1111111 : tail0=1'b0;
        16'b1110x0x0x1111111 : tail0=1'b0;
        16'b0x0x10x0x1111111 : tail0=1'b0;
        16'b110x10x0x1111111 : tail0=1'b0;
        16'b10x110x0x1111111 : tail0=1'b0;
        16'b0x1110x0x1111111 : tail0=1'b0;
        16'b111110x0x1111111 : tail0=1'b0;
        16'b0x0x0x10x1111111 : tail0=1'b0;
        16'b110x0x10x1111111 : tail0=1'b0;
        16'b10x10x10x1111111 : tail0=1'b0;
        16'b0x110x10x1111111 : tail0=1'b0;
        16'b11110x10x1111111 : tail0=1'b0;
        16'b10x0x110x1111111 : tail0=1'b0;
        16'b0x10x110x1111111 : tail0=1'b0;
        16'b1110x110x1111111 : tail0=1'b0;
        16'b0x0x1110x1111111 : tail0=1'b0;
        16'b110x1110x1111111 : tail0=1'b0;
        16'b10x11110x1111111 : tail0=1'b0;
        16'b0x111110x1111111 : tail0=1'b0;
        16'b11111110x1111111 : tail0=1'b0;
        16'b0x0x0x0x11111111 : tail0=1'b0;
        16'b110x0x0x11111111 : tail0=1'b0;
        16'b10x10x0x11111111 : tail0=1'b0;
        16'b0x110x0x11111111 : tail0=1'b0;
        16'b11110x0x11111111 : tail0=1'b0;
        16'b10x0x10x11111111 : tail0=1'b0;
        16'b0x10x10x11111111 : tail0=1'b0;
        16'b1110x10x11111111 : tail0=1'b0;
        16'b0x0x110x11111111 : tail0=1'b0;
        16'b110x110x11111111 : tail0=1'b0;
        16'b10x1110x11111111 : tail0=1'b0;
        16'b0x11110x11111111 : tail0=1'b0;
        16'b1111110x11111111 : tail0=1'b0;
        16'b10x0x0x111111111 : tail0=1'b0;
        16'b0x10x0x111111111 : tail0=1'b0;
        16'b1110x0x111111111 : tail0=1'b0;
        16'b0x0x10x111111111 : tail0=1'b0;
        16'b110x10x111111111 : tail0=1'b0;
        16'b10x110x111111111 : tail0=1'b0;
        16'b0x1110x111111111 : tail0=1'b0;
        16'b111110x111111111 : tail0=1'b0;
        16'b0x0x0x1111111111 : tail0=1'b0;
        16'b110x0x1111111111 : tail0=1'b0;
        16'b10x10x1111111111 : tail0=1'b0;
        16'b0x110x1111111111 : tail0=1'b0;
        16'b11110x1111111111 : tail0=1'b0;
        16'b10x0x11111111111 : tail0=1'b0;
        16'b0x10x11111111111 : tail0=1'b0;
        16'b1110x11111111111 : tail0=1'b0;
        16'b0x0x111111111111 : tail0=1'b0;
        16'b110x111111111111 : tail0=1'b0;
        16'b10x1111111111111 : tail0=1'b0;
        16'b0x11111111111111 : tail0=1'b0;
        16'b1111111111111111 : tail0=1'b0;
    endcase

  endfunction
