/*
Copyright 2022 Goran Dakov

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/


`define simd_padd 0
`define simd_psub 1
`define simd_paddsats 2
`define simd_psubsats 3
`define simd_paddsat 4
`define simd_psubsat 5
`define simd_pmins 6
`define simd_pmaxs 7
`define simd_pmin 8
`define simd_pmax 9
`define simd_cmp 10

`define simd_sar 11
`define simd_shr 12
`define simd_shl 13

`define simd_pand 16
`define simd_por 17
`define simd_pxor 18
`define simd_pmov 19
`define simd_pnand 20
`define simd_pnor 21
`define simd_pnxor 22
`define simd_pnot 23

