config.v