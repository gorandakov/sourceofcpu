`include "../struct.sv"

module fma_d(
  clk,
  rst,
  data_en,
  A,B,C,
  res,
  raise);
endmodule
