memop.v