/*
Copyright 2022 Goran Dakov

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

module frrv_rom(
  input [14:0] bits_in,
  output [14:0] bits_out);
  always @(bits_in) begin
    casex(bits_in)
        15'b0x0x0x0x0x0x0x0: bits_out=15'b010101010101010;
        15'b10x0x0x0x0x0x0x: bits_out=15'b101010101010101;
        15'b110x0x0x0x0x0x0: bits_out=15'b110101010101010;
        15'b0x10x0x0x0x0x0x: bits_out=15'b011010101010101;
        15'b1110x0x0x0x0x0x: bits_out=15'b111010101010101;
        15'b10x10x0x0x0x0x0: bits_out=15'b101101010101010;
        15'b0x110x0x0x0x0x0: bits_out=15'b011101010101010;
        15'b11110x0x0x0x0x0: bits_out=15'b111101010101010;
        15'b0x0x10x0x0x0x0x: bits_out=15'b010110101010101;
        15'b110x10x0x0x0x0x: bits_out=15'b110110101010101;
        15'b10x110x0x0x0x0x: bits_out=15'b101110101010101;
        15'b0x1110x0x0x0x0x: bits_out=15'b011110101010101;
        15'b111110x0x0x0x0x: bits_out=15'b111110101010101;
        15'b10x0x10x0x0x0x0: bits_out=15'b101011010101010;
        15'b0x10x10x0x0x0x0: bits_out=15'b011011010101010;
        15'b1110x10x0x0x0x0: bits_out=15'b111011010101010;
        15'b0x0x110x0x0x0x0: bits_out=15'b010111010101010;
        15'b110x110x0x0x0x0: bits_out=15'b110111010101010;
        15'b10x1110x0x0x0x0: bits_out=15'b101111010101010;
        15'b0x11110x0x0x0x0: bits_out=15'b011111010101010;
        15'b1111110x0x0x0x0: bits_out=15'b111111010101010;
        15'b0x0x0x10x0x0x0x: bits_out=15'b010101101010101;
        15'b110x0x10x0x0x0x: bits_out=15'b110101101010101;
        15'b10x10x10x0x0x0x: bits_out=15'b101101101010101;
        15'b0x110x10x0x0x0x: bits_out=15'b011101101010101;
        15'b11110x10x0x0x0x: bits_out=15'b111101101010101;
        15'b10x0x110x0x0x0x: bits_out=15'b101011101010101;
        15'b0x10x110x0x0x0x: bits_out=15'b011011101010101;
        15'b1110x110x0x0x0x: bits_out=15'b111011101010101;
        15'b0x0x1110x0x0x0x: bits_out=15'b010111101010101;
        15'b110x1110x0x0x0x: bits_out=15'b110111101010101;
        15'b10x11110x0x0x0x: bits_out=15'b101111101010101;
        15'b0x111110x0x0x0x: bits_out=15'b011111101010101;
        15'b11111110x0x0x0x: bits_out=15'b111111101010101;
        15'b10x0x0x10x0x0x0: bits_out=15'b101010110101010;
        15'b0x10x0x10x0x0x0: bits_out=15'b011010110101010;
        15'b1110x0x10x0x0x0: bits_out=15'b111010110101010;
        15'b0x0x10x10x0x0x0: bits_out=15'b010110110101010;
        15'b110x10x10x0x0x0: bits_out=15'b110110110101010;
        15'b10x110x10x0x0x0: bits_out=15'b101110110101010;
        15'b0x1110x10x0x0x0: bits_out=15'b011110110101010;
        15'b111110x10x0x0x0: bits_out=15'b111110110101010;
        15'b0x0x0x110x0x0x0: bits_out=15'b010101110101010;
        15'b110x0x110x0x0x0: bits_out=15'b110101110101010;
        15'b10x10x110x0x0x0: bits_out=15'b101101110101010;
        15'b0x110x110x0x0x0: bits_out=15'b011101110101010;
        15'b11110x110x0x0x0: bits_out=15'b111101110101010;
        15'b10x0x1110x0x0x0: bits_out=15'b101011110101010;
        15'b0x10x1110x0x0x0: bits_out=15'b011011110101010;
        15'b1110x1110x0x0x0: bits_out=15'b111011110101010;
        15'b0x0x11110x0x0x0: bits_out=15'b010111110101010;
        15'b110x11110x0x0x0: bits_out=15'b110111110101010;
        15'b10x111110x0x0x0: bits_out=15'b101111110101010;
        15'b0x1111110x0x0x0: bits_out=15'b011111110101010;
        15'b111111110x0x0x0: bits_out=15'b111111110101010;
        15'b0x0x0x0x10x0x0x: bits_out=15'b010101011010101;
        15'b110x0x0x10x0x0x: bits_out=15'b110101011010101;
        15'b10x10x0x10x0x0x: bits_out=15'b101101011010101;
        15'b0x110x0x10x0x0x: bits_out=15'b011101011010101;
        15'b11110x0x10x0x0x: bits_out=15'b111101011010101;
        15'b10x0x10x10x0x0x: bits_out=15'b101011011010101;
        15'b0x10x10x10x0x0x: bits_out=15'b011011011010101;
        15'b1110x10x10x0x0x: bits_out=15'b111011011010101;
        15'b0x0x110x10x0x0x: bits_out=15'b010111011010101;
        15'b110x110x10x0x0x: bits_out=15'b110111011010101;
        15'b10x1110x10x0x0x: bits_out=15'b101111011010101;
        15'b0x11110x10x0x0x: bits_out=15'b011111011010101;
        15'b1111110x10x0x0x: bits_out=15'b111111011010101;
        15'b10x0x0x110x0x0x: bits_out=15'b101010111010101;
        15'b0x10x0x110x0x0x: bits_out=15'b011010111010101;
        15'b1110x0x110x0x0x: bits_out=15'b111010111010101;
        15'b0x0x10x110x0x0x: bits_out=15'b010110111010101;
        15'b110x10x110x0x0x: bits_out=15'b110110111010101;
        15'b10x110x110x0x0x: bits_out=15'b101110111010101;
        15'b0x1110x110x0x0x: bits_out=15'b011110111010101;
        15'b111110x110x0x0x: bits_out=15'b111110111010101;
        15'b0x0x0x1110x0x0x: bits_out=15'b010101111010101;
        15'b110x0x1110x0x0x: bits_out=15'b110101111010101;
        15'b10x10x1110x0x0x: bits_out=15'b101101111010101;
        15'b0x110x1110x0x0x: bits_out=15'b011101111010101;
        15'b11110x1110x0x0x: bits_out=15'b111101111010101;
        15'b10x0x11110x0x0x: bits_out=15'b101011111010101;
        15'b0x10x11110x0x0x: bits_out=15'b011011111010101;
        15'b1110x11110x0x0x: bits_out=15'b111011111010101;
        15'b0x0x111110x0x0x: bits_out=15'b010111111010101;
        15'b110x111110x0x0x: bits_out=15'b110111111010101;
        15'b10x1111110x0x0x: bits_out=15'b101111111010101;
        15'b0x11111110x0x0x: bits_out=15'b011111111010101;
        15'b1111111110x0x0x: bits_out=15'b111111111010101;
        15'b10x0x0x0x10x0x0: bits_out=15'b101010101101010;
        15'b0x10x0x0x10x0x0: bits_out=15'b011010101101010;
        15'b1110x0x0x10x0x0: bits_out=15'b111010101101010;
        15'b0x0x10x0x10x0x0: bits_out=15'b010110101101010;
        15'b110x10x0x10x0x0: bits_out=15'b110110101101010;
        15'b10x110x0x10x0x0: bits_out=15'b101110101101010;
        15'b0x1110x0x10x0x0: bits_out=15'b011110101101010;
        15'b111110x0x10x0x0: bits_out=15'b111110101101010;
        15'b0x0x0x10x10x0x0: bits_out=15'b010101101101010;
        15'b110x0x10x10x0x0: bits_out=15'b110101101101010;
        15'b10x10x10x10x0x0: bits_out=15'b101101101101010;
        15'b0x110x10x10x0x0: bits_out=15'b011101101101010;
        15'b11110x10x10x0x0: bits_out=15'b111101101101010;
        15'b10x0x110x10x0x0: bits_out=15'b101011101101010;
        15'b0x10x110x10x0x0: bits_out=15'b011011101101010;
        15'b1110x110x10x0x0: bits_out=15'b111011101101010;
        15'b0x0x1110x10x0x0: bits_out=15'b010111101101010;
        15'b110x1110x10x0x0: bits_out=15'b110111101101010;
        15'b10x11110x10x0x0: bits_out=15'b101111101101010;
        15'b0x111110x10x0x0: bits_out=15'b011111101101010;
        15'b11111110x10x0x0: bits_out=15'b111111101101010;
        15'b0x0x0x0x110x0x0: bits_out=15'b010101011101010;
        15'b110x0x0x110x0x0: bits_out=15'b110101011101010;
        15'b10x10x0x110x0x0: bits_out=15'b101101011101010;
        15'b0x110x0x110x0x0: bits_out=15'b011101011101010;
        15'b11110x0x110x0x0: bits_out=15'b111101011101010;
        15'b10x0x10x110x0x0: bits_out=15'b101011011101010;
        15'b0x10x10x110x0x0: bits_out=15'b011011011101010;
        15'b1110x10x110x0x0: bits_out=15'b111011011101010;
        15'b0x0x110x110x0x0: bits_out=15'b010111011101010;
        15'b110x110x110x0x0: bits_out=15'b110111011101010;
        15'b10x1110x110x0x0: bits_out=15'b101111011101010;
        15'b0x11110x110x0x0: bits_out=15'b011111011101010;
        15'b1111110x110x0x0: bits_out=15'b111111011101010;
        15'b10x0x0x1110x0x0: bits_out=15'b101010111101010;
        15'b0x10x0x1110x0x0: bits_out=15'b011010111101010;
        15'b1110x0x1110x0x0: bits_out=15'b111010111101010;
        15'b0x0x10x1110x0x0: bits_out=15'b010110111101010;
        15'b110x10x1110x0x0: bits_out=15'b110110111101010;
        15'b10x110x1110x0x0: bits_out=15'b101110111101010;
        15'b0x1110x1110x0x0: bits_out=15'b011110111101010;
        15'b111110x1110x0x0: bits_out=15'b111110111101010;
        15'b0x0x0x11110x0x0: bits_out=15'b010101111101010;
        15'b110x0x11110x0x0: bits_out=15'b110101111101010;
        15'b10x10x11110x0x0: bits_out=15'b101101111101010;
        15'b0x110x11110x0x0: bits_out=15'b011101111101010;
        15'b11110x11110x0x0: bits_out=15'b111101111101010;
        15'b10x0x111110x0x0: bits_out=15'b101011111101010;
        15'b0x10x111110x0x0: bits_out=15'b011011111101010;
        15'b1110x111110x0x0: bits_out=15'b111011111101010;
        15'b0x0x1111110x0x0: bits_out=15'b010111111101010;
        15'b110x1111110x0x0: bits_out=15'b110111111101010;
        15'b10x11111110x0x0: bits_out=15'b101111111101010;
        15'b0x111111110x0x0: bits_out=15'b011111111101010;
        15'b11111111110x0x0: bits_out=15'b111111111101010;
        15'b0x0x0x0x0x10x0x: bits_out=15'b010101010110101;
        15'b110x0x0x0x10x0x: bits_out=15'b110101010110101;
        15'b10x10x0x0x10x0x: bits_out=15'b101101010110101;
        15'b0x110x0x0x10x0x: bits_out=15'b011101010110101;
        15'b11110x0x0x10x0x: bits_out=15'b111101010110101;
        15'b10x0x10x0x10x0x: bits_out=15'b101011010110101;
        15'b0x10x10x0x10x0x: bits_out=15'b011011010110101;
        15'b1110x10x0x10x0x: bits_out=15'b111011010110101;
        15'b0x0x110x0x10x0x: bits_out=15'b010111010110101;
        15'b110x110x0x10x0x: bits_out=15'b110111010110101;
        15'b10x1110x0x10x0x: bits_out=15'b101111010110101;
        15'b0x11110x0x10x0x: bits_out=15'b011111010110101;
        15'b1111110x0x10x0x: bits_out=15'b111111010110101;
        15'b10x0x0x10x10x0x: bits_out=15'b101010110110101;
        15'b0x10x0x10x10x0x: bits_out=15'b011010110110101;
        15'b1110x0x10x10x0x: bits_out=15'b111010110110101;
        15'b0x0x10x10x10x0x: bits_out=15'b010110110110101;
        15'b110x10x10x10x0x: bits_out=15'b110110110110101;
        15'b10x110x10x10x0x: bits_out=15'b101110110110101;
        15'b0x1110x10x10x0x: bits_out=15'b011110110110101;
        15'b111110x10x10x0x: bits_out=15'b111110110110101;
        15'b0x0x0x110x10x0x: bits_out=15'b010101110110101;
        15'b110x0x110x10x0x: bits_out=15'b110101110110101;
        15'b10x10x110x10x0x: bits_out=15'b101101110110101;
        15'b0x110x110x10x0x: bits_out=15'b011101110110101;
        15'b11110x110x10x0x: bits_out=15'b111101110110101;
        15'b10x0x1110x10x0x: bits_out=15'b101011110110101;
        15'b0x10x1110x10x0x: bits_out=15'b011011110110101;
        15'b1110x1110x10x0x: bits_out=15'b111011110110101;
        15'b0x0x11110x10x0x: bits_out=15'b010111110110101;
        15'b110x11110x10x0x: bits_out=15'b110111110110101;
        15'b10x111110x10x0x: bits_out=15'b101111110110101;
        15'b0x1111110x10x0x: bits_out=15'b011111110110101;
        15'b111111110x10x0x: bits_out=15'b111111110110101;
        15'b10x0x0x0x110x0x: bits_out=15'b101010101110101;
        15'b0x10x0x0x110x0x: bits_out=15'b011010101110101;
        15'b1110x0x0x110x0x: bits_out=15'b111010101110101;
        15'b0x0x10x0x110x0x: bits_out=15'b010110101110101;
        15'b110x10x0x110x0x: bits_out=15'b110110101110101;
        15'b10x110x0x110x0x: bits_out=15'b101110101110101;
        15'b0x1110x0x110x0x: bits_out=15'b011110101110101;
        15'b111110x0x110x0x: bits_out=15'b111110101110101;
        15'b0x0x0x10x110x0x: bits_out=15'b010101101110101;
        15'b110x0x10x110x0x: bits_out=15'b110101101110101;
        15'b10x10x10x110x0x: bits_out=15'b101101101110101;
        15'b0x110x10x110x0x: bits_out=15'b011101101110101;
        15'b11110x10x110x0x: bits_out=15'b111101101110101;
        15'b10x0x110x110x0x: bits_out=15'b101011101110101;
        15'b0x10x110x110x0x: bits_out=15'b011011101110101;
        15'b1110x110x110x0x: bits_out=15'b111011101110101;
        15'b0x0x1110x110x0x: bits_out=15'b010111101110101;
        15'b110x1110x110x0x: bits_out=15'b110111101110101;
        15'b10x11110x110x0x: bits_out=15'b101111101110101;
        15'b0x111110x110x0x: bits_out=15'b011111101110101;
        15'b11111110x110x0x: bits_out=15'b111111101110101;
        15'b0x0x0x0x1110x0x: bits_out=15'b010101011110101;
        15'b110x0x0x1110x0x: bits_out=15'b110101011110101;
        15'b10x10x0x1110x0x: bits_out=15'b101101011110101;
        15'b0x110x0x1110x0x: bits_out=15'b011101011110101;
        15'b11110x0x1110x0x: bits_out=15'b111101011110101;
        15'b10x0x10x1110x0x: bits_out=15'b101011011110101;
        15'b0x10x10x1110x0x: bits_out=15'b011011011110101;
        15'b1110x10x1110x0x: bits_out=15'b111011011110101;
        15'b0x0x110x1110x0x: bits_out=15'b010111011110101;
        15'b110x110x1110x0x: bits_out=15'b110111011110101;
        15'b10x1110x1110x0x: bits_out=15'b101111011110101;
        15'b0x11110x1110x0x: bits_out=15'b011111011110101;
        15'b1111110x1110x0x: bits_out=15'b111111011110101;
        15'b10x0x0x11110x0x: bits_out=15'b101010111110101;
        15'b0x10x0x11110x0x: bits_out=15'b011010111110101;
        15'b1110x0x11110x0x: bits_out=15'b111010111110101;
        15'b0x0x10x11110x0x: bits_out=15'b010110111110101;
        15'b110x10x11110x0x: bits_out=15'b110110111110101;
        15'b10x110x11110x0x: bits_out=15'b101110111110101;
        15'b0x1110x11110x0x: bits_out=15'b011110111110101;
        15'b111110x11110x0x: bits_out=15'b111110111110101;
        15'b0x0x0x111110x0x: bits_out=15'b010101111110101;
        15'b110x0x111110x0x: bits_out=15'b110101111110101;
        15'b10x10x111110x0x: bits_out=15'b101101111110101;
        15'b0x110x111110x0x: bits_out=15'b011101111110101;
        15'b11110x111110x0x: bits_out=15'b111101111110101;
        15'b10x0x1111110x0x: bits_out=15'b101011111110101;
        15'b0x10x1111110x0x: bits_out=15'b011011111110101;
        15'b1110x1111110x0x: bits_out=15'b111011111110101;
        15'b0x0x11111110x0x: bits_out=15'b010111111110101;
        15'b110x11111110x0x: bits_out=15'b110111111110101;
        15'b10x111111110x0x: bits_out=15'b101111111110101;
        15'b0x1111111110x0x: bits_out=15'b011111111110101;
        15'b111111111110x0x: bits_out=15'b111111111110101;
        15'b10x0x0x0x0x10x0: bits_out=15'b101010101011010;
        15'b0x10x0x0x0x10x0: bits_out=15'b011010101011010;
        15'b1110x0x0x0x10x0: bits_out=15'b111010101011010;
        15'b0x0x10x0x0x10x0: bits_out=15'b010110101011010;
        15'b110x10x0x0x10x0: bits_out=15'b110110101011010;
        15'b10x110x0x0x10x0: bits_out=15'b101110101011010;
        15'b0x1110x0x0x10x0: bits_out=15'b011110101011010;
        15'b111110x0x0x10x0: bits_out=15'b111110101011010;
        15'b0x0x0x10x0x10x0: bits_out=15'b010101101011010;
        15'b110x0x10x0x10x0: bits_out=15'b110101101011010;
        15'b10x10x10x0x10x0: bits_out=15'b101101101011010;
        15'b0x110x10x0x10x0: bits_out=15'b011101101011010;
        15'b11110x10x0x10x0: bits_out=15'b111101101011010;
        15'b10x0x110x0x10x0: bits_out=15'b101011101011010;
        15'b0x10x110x0x10x0: bits_out=15'b011011101011010;
        15'b1110x110x0x10x0: bits_out=15'b111011101011010;
        15'b0x0x1110x0x10x0: bits_out=15'b010111101011010;
        15'b110x1110x0x10x0: bits_out=15'b110111101011010;
        15'b10x11110x0x10x0: bits_out=15'b101111101011010;
        15'b0x111110x0x10x0: bits_out=15'b011111101011010;
        15'b11111110x0x10x0: bits_out=15'b111111101011010;
        15'b0x0x0x0x10x10x0: bits_out=15'b010101011011010;
        15'b110x0x0x10x10x0: bits_out=15'b110101011011010;
        15'b10x10x0x10x10x0: bits_out=15'b101101011011010;
        15'b0x110x0x10x10x0: bits_out=15'b011101011011010;
        15'b11110x0x10x10x0: bits_out=15'b111101011011010;
        15'b10x0x10x10x10x0: bits_out=15'b101011011011010;
        15'b0x10x10x10x10x0: bits_out=15'b011011011011010;
        15'b1110x10x10x10x0: bits_out=15'b111011011011010;
        15'b0x0x110x10x10x0: bits_out=15'b010111011011010;
        15'b110x110x10x10x0: bits_out=15'b110111011011010;
        15'b10x1110x10x10x0: bits_out=15'b101111011011010;
        15'b0x11110x10x10x0: bits_out=15'b011111011011010;
        15'b1111110x10x10x0: bits_out=15'b111111011011010;
        15'b10x0x0x110x10x0: bits_out=15'b101010111011010;
        15'b0x10x0x110x10x0: bits_out=15'b011010111011010;
        15'b1110x0x110x10x0: bits_out=15'b111010111011010;
        15'b0x0x10x110x10x0: bits_out=15'b010110111011010;
        15'b110x10x110x10x0: bits_out=15'b110110111011010;
        15'b10x110x110x10x0: bits_out=15'b101110111011010;
        15'b0x1110x110x10x0: bits_out=15'b011110111011010;
        15'b111110x110x10x0: bits_out=15'b111110111011010;
        15'b0x0x0x1110x10x0: bits_out=15'b010101111011010;
        15'b110x0x1110x10x0: bits_out=15'b110101111011010;
        15'b10x10x1110x10x0: bits_out=15'b101101111011010;
        15'b0x110x1110x10x0: bits_out=15'b011101111011010;
        15'b11110x1110x10x0: bits_out=15'b111101111011010;
        15'b10x0x11110x10x0: bits_out=15'b101011111011010;
        15'b0x10x11110x10x0: bits_out=15'b011011111011010;
        15'b1110x11110x10x0: bits_out=15'b111011111011010;
        15'b0x0x111110x10x0: bits_out=15'b010111111011010;
        15'b110x111110x10x0: bits_out=15'b110111111011010;
        15'b10x1111110x10x0: bits_out=15'b101111111011010;
        15'b0x11111110x10x0: bits_out=15'b011111111011010;
        15'b1111111110x10x0: bits_out=15'b111111111011010;
        15'b0x0x0x0x0x110x0: bits_out=15'b010101010111010;
        15'b110x0x0x0x110x0: bits_out=15'b110101010111010;
        15'b10x10x0x0x110x0: bits_out=15'b101101010111010;
        15'b0x110x0x0x110x0: bits_out=15'b011101010111010;
        15'b11110x0x0x110x0: bits_out=15'b111101010111010;
        15'b10x0x10x0x110x0: bits_out=15'b101011010111010;
        15'b0x10x10x0x110x0: bits_out=15'b011011010111010;
        15'b1110x10x0x110x0: bits_out=15'b111011010111010;
        15'b0x0x110x0x110x0: bits_out=15'b010111010111010;
        15'b110x110x0x110x0: bits_out=15'b110111010111010;
        15'b10x1110x0x110x0: bits_out=15'b101111010111010;
        15'b0x11110x0x110x0: bits_out=15'b011111010111010;
        15'b1111110x0x110x0: bits_out=15'b111111010111010;
        15'b10x0x0x10x110x0: bits_out=15'b101010110111010;
        15'b0x10x0x10x110x0: bits_out=15'b011010110111010;
        15'b1110x0x10x110x0: bits_out=15'b111010110111010;
        15'b0x0x10x10x110x0: bits_out=15'b010110110111010;
        15'b110x10x10x110x0: bits_out=15'b110110110111010;
        15'b10x110x10x110x0: bits_out=15'b101110110111010;
        15'b0x1110x10x110x0: bits_out=15'b011110110111010;
        15'b111110x10x110x0: bits_out=15'b111110110111010;
        15'b0x0x0x110x110x0: bits_out=15'b010101110111010;
        15'b110x0x110x110x0: bits_out=15'b110101110111010;
        15'b10x10x110x110x0: bits_out=15'b101101110111010;
        15'b0x110x110x110x0: bits_out=15'b011101110111010;
        15'b11110x110x110x0: bits_out=15'b111101110111010;
        15'b10x0x1110x110x0: bits_out=15'b101011110111010;
        15'b0x10x1110x110x0: bits_out=15'b011011110111010;
        15'b1110x1110x110x0: bits_out=15'b111011110111010;
        15'b0x0x11110x110x0: bits_out=15'b010111110111010;
        15'b110x11110x110x0: bits_out=15'b110111110111010;
        15'b10x111110x110x0: bits_out=15'b101111110111010;
        15'b0x1111110x110x0: bits_out=15'b011111110111010;
        15'b111111110x110x0: bits_out=15'b111111110111010;
        15'b10x0x0x0x1110x0: bits_out=15'b101010101111010;
        15'b0x10x0x0x1110x0: bits_out=15'b011010101111010;
        15'b1110x0x0x1110x0: bits_out=15'b111010101111010;
        15'b0x0x10x0x1110x0: bits_out=15'b010110101111010;
        15'b110x10x0x1110x0: bits_out=15'b110110101111010;
        15'b10x110x0x1110x0: bits_out=15'b101110101111010;
        15'b0x1110x0x1110x0: bits_out=15'b011110101111010;
        15'b111110x0x1110x0: bits_out=15'b111110101111010;
        15'b0x0x0x10x1110x0: bits_out=15'b010101101111010;
        15'b110x0x10x1110x0: bits_out=15'b110101101111010;
        15'b10x10x10x1110x0: bits_out=15'b101101101111010;
        15'b0x110x10x1110x0: bits_out=15'b011101101111010;
        15'b11110x10x1110x0: bits_out=15'b111101101111010;
        15'b10x0x110x1110x0: bits_out=15'b101011101111010;
        15'b0x10x110x1110x0: bits_out=15'b011011101111010;
        15'b1110x110x1110x0: bits_out=15'b111011101111010;
        15'b0x0x1110x1110x0: bits_out=15'b010111101111010;
        15'b110x1110x1110x0: bits_out=15'b110111101111010;
        15'b10x11110x1110x0: bits_out=15'b101111101111010;
        15'b0x111110x1110x0: bits_out=15'b011111101111010;
        15'b11111110x1110x0: bits_out=15'b111111101111010;
        15'b0x0x0x0x11110x0: bits_out=15'b010101011111010;
        15'b110x0x0x11110x0: bits_out=15'b110101011111010;
        15'b10x10x0x11110x0: bits_out=15'b101101011111010;
        15'b0x110x0x11110x0: bits_out=15'b011101011111010;
        15'b11110x0x11110x0: bits_out=15'b111101011111010;
        15'b10x0x10x11110x0: bits_out=15'b101011011111010;
        15'b0x10x10x11110x0: bits_out=15'b011011011111010;
        15'b1110x10x11110x0: bits_out=15'b111011011111010;
        15'b0x0x110x11110x0: bits_out=15'b010111011111010;
        15'b110x110x11110x0: bits_out=15'b110111011111010;
        15'b10x1110x11110x0: bits_out=15'b101111011111010;
        15'b0x11110x11110x0: bits_out=15'b011111011111010;
        15'b1111110x11110x0: bits_out=15'b111111011111010;
        15'b10x0x0x111110x0: bits_out=15'b101010111111010;
        15'b0x10x0x111110x0: bits_out=15'b011010111111010;
        15'b1110x0x111110x0: bits_out=15'b111010111111010;
        15'b0x0x10x111110x0: bits_out=15'b010110111111010;
        15'b110x10x111110x0: bits_out=15'b110110111111010;
        15'b10x110x111110x0: bits_out=15'b101110111111010;
        15'b0x1110x111110x0: bits_out=15'b011110111111010;
        15'b111110x111110x0: bits_out=15'b111110111111010;
        15'b0x0x0x1111110x0: bits_out=15'b010101111111010;
        15'b110x0x1111110x0: bits_out=15'b110101111111010;
        15'b10x10x1111110x0: bits_out=15'b101101111111010;
        15'b0x110x1111110x0: bits_out=15'b011101111111010;
        15'b11110x1111110x0: bits_out=15'b111101111111010;
        15'b10x0x11111110x0: bits_out=15'b101011111111010;
        15'b0x10x11111110x0: bits_out=15'b011011111111010;
        15'b1110x11111110x0: bits_out=15'b111011111111010;
        15'b0x0x111111110x0: bits_out=15'b010111111111010;
        15'b110x111111110x0: bits_out=15'b110111111111010;
        15'b10x1111111110x0: bits_out=15'b101111111111010;
        15'b0x11111111110x0: bits_out=15'b011111111111010;
        15'b1111111111110x0: bits_out=15'b111111111111010;
        15'b0x0x0x0x0x0x10x: bits_out=15'b010101010101101;
        15'b110x0x0x0x0x10x: bits_out=15'b110101010101101;
        15'b10x10x0x0x0x10x: bits_out=15'b101101010101101;
        15'b0x110x0x0x0x10x: bits_out=15'b011101010101101;
        15'b11110x0x0x0x10x: bits_out=15'b111101010101101;
        15'b10x0x10x0x0x10x: bits_out=15'b101011010101101;
        15'b0x10x10x0x0x10x: bits_out=15'b011011010101101;
        15'b1110x10x0x0x10x: bits_out=15'b111011010101101;
        15'b0x0x110x0x0x10x: bits_out=15'b010111010101101;
        15'b110x110x0x0x10x: bits_out=15'b110111010101101;
        15'b10x1110x0x0x10x: bits_out=15'b101111010101101;
        15'b0x11110x0x0x10x: bits_out=15'b011111010101101;
        15'b1111110x0x0x10x: bits_out=15'b111111010101101;
        15'b10x0x0x10x0x10x: bits_out=15'b101010110101101;
        15'b0x10x0x10x0x10x: bits_out=15'b011010110101101;
        15'b1110x0x10x0x10x: bits_out=15'b111010110101101;
        15'b0x0x10x10x0x10x: bits_out=15'b010110110101101;
        15'b110x10x10x0x10x: bits_out=15'b110110110101101;
        15'b10x110x10x0x10x: bits_out=15'b101110110101101;
        15'b0x1110x10x0x10x: bits_out=15'b011110110101101;
        15'b111110x10x0x10x: bits_out=15'b111110110101101;
        15'b0x0x0x110x0x10x: bits_out=15'b010101110101101;
        15'b110x0x110x0x10x: bits_out=15'b110101110101101;
        15'b10x10x110x0x10x: bits_out=15'b101101110101101;
        15'b0x110x110x0x10x: bits_out=15'b011101110101101;
        15'b11110x110x0x10x: bits_out=15'b111101110101101;
        15'b10x0x1110x0x10x: bits_out=15'b101011110101101;
        15'b0x10x1110x0x10x: bits_out=15'b011011110101101;
        15'b1110x1110x0x10x: bits_out=15'b111011110101101;
        15'b0x0x11110x0x10x: bits_out=15'b010111110101101;
        15'b110x11110x0x10x: bits_out=15'b110111110101101;
        15'b10x111110x0x10x: bits_out=15'b101111110101101;
        15'b0x1111110x0x10x: bits_out=15'b011111110101101;
        15'b111111110x0x10x: bits_out=15'b111111110101101;
        15'b10x0x0x0x10x10x: bits_out=15'b101010101101101;
        15'b0x10x0x0x10x10x: bits_out=15'b011010101101101;
        15'b1110x0x0x10x10x: bits_out=15'b111010101101101;
        15'b0x0x10x0x10x10x: bits_out=15'b010110101101101;
        15'b110x10x0x10x10x: bits_out=15'b110110101101101;
        15'b10x110x0x10x10x: bits_out=15'b101110101101101;
        15'b0x1110x0x10x10x: bits_out=15'b011110101101101;
        15'b111110x0x10x10x: bits_out=15'b111110101101101;
        15'b0x0x0x10x10x10x: bits_out=15'b010101101101101;
        15'b110x0x10x10x10x: bits_out=15'b110101101101101;
        15'b10x10x10x10x10x: bits_out=15'b101101101101101;
        15'b0x110x10x10x10x: bits_out=15'b011101101101101;
        15'b11110x10x10x10x: bits_out=15'b111101101101101;
        15'b10x0x110x10x10x: bits_out=15'b101011101101101;
        15'b0x10x110x10x10x: bits_out=15'b011011101101101;
        15'b1110x110x10x10x: bits_out=15'b111011101101101;
        15'b0x0x1110x10x10x: bits_out=15'b010111101101101;
        15'b110x1110x10x10x: bits_out=15'b110111101101101;
        15'b10x11110x10x10x: bits_out=15'b101111101101101;
        15'b0x111110x10x10x: bits_out=15'b011111101101101;
        15'b11111110x10x10x: bits_out=15'b111111101101101;
        15'b0x0x0x0x110x10x: bits_out=15'b010101011101101;
        15'b110x0x0x110x10x: bits_out=15'b110101011101101;
        15'b10x10x0x110x10x: bits_out=15'b101101011101101;
        15'b0x110x0x110x10x: bits_out=15'b011101011101101;
        15'b11110x0x110x10x: bits_out=15'b111101011101101;
        15'b10x0x10x110x10x: bits_out=15'b101011011101101;
        15'b0x10x10x110x10x: bits_out=15'b011011011101101;
        15'b1110x10x110x10x: bits_out=15'b111011011101101;
        15'b0x0x110x110x10x: bits_out=15'b010111011101101;
        15'b110x110x110x10x: bits_out=15'b110111011101101;
        15'b10x1110x110x10x: bits_out=15'b101111011101101;
        15'b0x11110x110x10x: bits_out=15'b011111011101101;
        15'b1111110x110x10x: bits_out=15'b111111011101101;
        15'b10x0x0x1110x10x: bits_out=15'b101010111101101;
        15'b0x10x0x1110x10x: bits_out=15'b011010111101101;
        15'b1110x0x1110x10x: bits_out=15'b111010111101101;
        15'b0x0x10x1110x10x: bits_out=15'b010110111101101;
        15'b110x10x1110x10x: bits_out=15'b110110111101101;
        15'b10x110x1110x10x: bits_out=15'b101110111101101;
        15'b0x1110x1110x10x: bits_out=15'b011110111101101;
        15'b111110x1110x10x: bits_out=15'b111110111101101;
        15'b0x0x0x11110x10x: bits_out=15'b010101111101101;
        15'b110x0x11110x10x: bits_out=15'b110101111101101;
        15'b10x10x11110x10x: bits_out=15'b101101111101101;
        15'b0x110x11110x10x: bits_out=15'b011101111101101;
        15'b11110x11110x10x: bits_out=15'b111101111101101;
        15'b10x0x111110x10x: bits_out=15'b101011111101101;
        15'b0x10x111110x10x: bits_out=15'b011011111101101;
        15'b1110x111110x10x: bits_out=15'b111011111101101;
        15'b0x0x1111110x10x: bits_out=15'b010111111101101;
        15'b110x1111110x10x: bits_out=15'b110111111101101;
        15'b10x11111110x10x: bits_out=15'b101111111101101;
        15'b0x111111110x10x: bits_out=15'b011111111101101;
        15'b11111111110x10x: bits_out=15'b111111111101101;
        15'b10x0x0x0x0x110x: bits_out=15'b101010101011101;
        15'b0x10x0x0x0x110x: bits_out=15'b011010101011101;
        15'b1110x0x0x0x110x: bits_out=15'b111010101011101;
        15'b0x0x10x0x0x110x: bits_out=15'b010110101011101;
        15'b110x10x0x0x110x: bits_out=15'b110110101011101;
        15'b10x110x0x0x110x: bits_out=15'b101110101011101;
        15'b0x1110x0x0x110x: bits_out=15'b011110101011101;
        15'b111110x0x0x110x: bits_out=15'b111110101011101;
        15'b0x0x0x10x0x110x: bits_out=15'b010101101011101;
        15'b110x0x10x0x110x: bits_out=15'b110101101011101;
        15'b10x10x10x0x110x: bits_out=15'b101101101011101;
        15'b0x110x10x0x110x: bits_out=15'b011101101011101;
        15'b11110x10x0x110x: bits_out=15'b111101101011101;
        15'b10x0x110x0x110x: bits_out=15'b101011101011101;
        15'b0x10x110x0x110x: bits_out=15'b011011101011101;
        15'b1110x110x0x110x: bits_out=15'b111011101011101;
        15'b0x0x1110x0x110x: bits_out=15'b010111101011101;
        15'b110x1110x0x110x: bits_out=15'b110111101011101;
        15'b10x11110x0x110x: bits_out=15'b101111101011101;
        15'b0x111110x0x110x: bits_out=15'b011111101011101;
        15'b11111110x0x110x: bits_out=15'b111111101011101;
        15'b0x0x0x0x10x110x: bits_out=15'b010101011011101;
        15'b110x0x0x10x110x: bits_out=15'b110101011011101;
        15'b10x10x0x10x110x: bits_out=15'b101101011011101;
        15'b0x110x0x10x110x: bits_out=15'b011101011011101;
        15'b11110x0x10x110x: bits_out=15'b111101011011101;
        15'b10x0x10x10x110x: bits_out=15'b101011011011101;
        15'b0x10x10x10x110x: bits_out=15'b011011011011101;
        15'b1110x10x10x110x: bits_out=15'b111011011011101;
        15'b0x0x110x10x110x: bits_out=15'b010111011011101;
        15'b110x110x10x110x: bits_out=15'b110111011011101;
        15'b10x1110x10x110x: bits_out=15'b101111011011101;
        15'b0x11110x10x110x: bits_out=15'b011111011011101;
        15'b1111110x10x110x: bits_out=15'b111111011011101;
        15'b10x0x0x110x110x: bits_out=15'b101010111011101;
        15'b0x10x0x110x110x: bits_out=15'b011010111011101;
        15'b1110x0x110x110x: bits_out=15'b111010111011101;
        15'b0x0x10x110x110x: bits_out=15'b010110111011101;
        15'b110x10x110x110x: bits_out=15'b110110111011101;
        15'b10x110x110x110x: bits_out=15'b101110111011101;
        15'b0x1110x110x110x: bits_out=15'b011110111011101;
        15'b111110x110x110x: bits_out=15'b111110111011101;
        15'b0x0x0x1110x110x: bits_out=15'b010101111011101;
        15'b110x0x1110x110x: bits_out=15'b110101111011101;
        15'b10x10x1110x110x: bits_out=15'b101101111011101;
        15'b0x110x1110x110x: bits_out=15'b011101111011101;
        15'b11110x1110x110x: bits_out=15'b111101111011101;
        15'b10x0x11110x110x: bits_out=15'b101011111011101;
        15'b0x10x11110x110x: bits_out=15'b011011111011101;
        15'b1110x11110x110x: bits_out=15'b111011111011101;
        15'b0x0x111110x110x: bits_out=15'b010111111011101;
        15'b110x111110x110x: bits_out=15'b110111111011101;
        15'b10x1111110x110x: bits_out=15'b101111111011101;
        15'b0x11111110x110x: bits_out=15'b011111111011101;
        15'b1111111110x110x: bits_out=15'b111111111011101;
        15'b0x0x0x0x0x1110x: bits_out=15'b010101010111101;
        15'b110x0x0x0x1110x: bits_out=15'b110101010111101;
        15'b10x10x0x0x1110x: bits_out=15'b101101010111101;
        15'b0x110x0x0x1110x: bits_out=15'b011101010111101;
        15'b11110x0x0x1110x: bits_out=15'b111101010111101;
        15'b10x0x10x0x1110x: bits_out=15'b101011010111101;
        15'b0x10x10x0x1110x: bits_out=15'b011011010111101;
        15'b1110x10x0x1110x: bits_out=15'b111011010111101;
        15'b0x0x110x0x1110x: bits_out=15'b010111010111101;
        15'b110x110x0x1110x: bits_out=15'b110111010111101;
        15'b10x1110x0x1110x: bits_out=15'b101111010111101;
        15'b0x11110x0x1110x: bits_out=15'b011111010111101;
        15'b1111110x0x1110x: bits_out=15'b111111010111101;
        15'b10x0x0x10x1110x: bits_out=15'b101010110111101;
        15'b0x10x0x10x1110x: bits_out=15'b011010110111101;
        15'b1110x0x10x1110x: bits_out=15'b111010110111101;
        15'b0x0x10x10x1110x: bits_out=15'b010110110111101;
        15'b110x10x10x1110x: bits_out=15'b110110110111101;
        15'b10x110x10x1110x: bits_out=15'b101110110111101;
        15'b0x1110x10x1110x: bits_out=15'b011110110111101;
        15'b111110x10x1110x: bits_out=15'b111110110111101;
        15'b0x0x0x110x1110x: bits_out=15'b010101110111101;
        15'b110x0x110x1110x: bits_out=15'b110101110111101;
        15'b10x10x110x1110x: bits_out=15'b101101110111101;
        15'b0x110x110x1110x: bits_out=15'b011101110111101;
        15'b11110x110x1110x: bits_out=15'b111101110111101;
        15'b10x0x1110x1110x: bits_out=15'b101011110111101;
        15'b0x10x1110x1110x: bits_out=15'b011011110111101;
        15'b1110x1110x1110x: bits_out=15'b111011110111101;
        15'b0x0x11110x1110x: bits_out=15'b010111110111101;
        15'b110x11110x1110x: bits_out=15'b110111110111101;
        15'b10x111110x1110x: bits_out=15'b101111110111101;
        15'b0x1111110x1110x: bits_out=15'b011111110111101;
        15'b111111110x1110x: bits_out=15'b111111110111101;
        15'b10x0x0x0x11110x: bits_out=15'b101010101111101;
        15'b0x10x0x0x11110x: bits_out=15'b011010101111101;
        15'b1110x0x0x11110x: bits_out=15'b111010101111101;
        15'b0x0x10x0x11110x: bits_out=15'b010110101111101;
        15'b110x10x0x11110x: bits_out=15'b110110101111101;
        15'b10x110x0x11110x: bits_out=15'b101110101111101;
        15'b0x1110x0x11110x: bits_out=15'b011110101111101;
        15'b111110x0x11110x: bits_out=15'b111110101111101;
        15'b0x0x0x10x11110x: bits_out=15'b010101101111101;
        15'b110x0x10x11110x: bits_out=15'b110101101111101;
        15'b10x10x10x11110x: bits_out=15'b101101101111101;
        15'b0x110x10x11110x: bits_out=15'b011101101111101;
        15'b11110x10x11110x: bits_out=15'b111101101111101;
        15'b10x0x110x11110x: bits_out=15'b101011101111101;
        15'b0x10x110x11110x: bits_out=15'b011011101111101;
        15'b1110x110x11110x: bits_out=15'b111011101111101;
        15'b0x0x1110x11110x: bits_out=15'b010111101111101;
        15'b110x1110x11110x: bits_out=15'b110111101111101;
        15'b10x11110x11110x: bits_out=15'b101111101111101;
        15'b0x111110x11110x: bits_out=15'b011111101111101;
        15'b11111110x11110x: bits_out=15'b111111101111101;
        15'b0x0x0x0x111110x: bits_out=15'b010101011111101;
        15'b110x0x0x111110x: bits_out=15'b110101011111101;
        15'b10x10x0x111110x: bits_out=15'b101101011111101;
        15'b0x110x0x111110x: bits_out=15'b011101011111101;
        15'b11110x0x111110x: bits_out=15'b111101011111101;
        15'b10x0x10x111110x: bits_out=15'b101011011111101;
        15'b0x10x10x111110x: bits_out=15'b011011011111101;
        15'b1110x10x111110x: bits_out=15'b111011011111101;
        15'b0x0x110x111110x: bits_out=15'b010111011111101;
        15'b110x110x111110x: bits_out=15'b110111011111101;
        15'b10x1110x111110x: bits_out=15'b101111011111101;
        15'b0x11110x111110x: bits_out=15'b011111011111101;
        15'b1111110x111110x: bits_out=15'b111111011111101;
        15'b10x0x0x1111110x: bits_out=15'b101010111111101;
        15'b0x10x0x1111110x: bits_out=15'b011010111111101;
        15'b1110x0x1111110x: bits_out=15'b111010111111101;
        15'b0x0x10x1111110x: bits_out=15'b010110111111101;
        15'b110x10x1111110x: bits_out=15'b110110111111101;
        15'b10x110x1111110x: bits_out=15'b101110111111101;
        15'b0x1110x1111110x: bits_out=15'b011110111111101;
        15'b111110x1111110x: bits_out=15'b111110111111101;
        15'b0x0x0x11111110x: bits_out=15'b010101111111101;
        15'b110x0x11111110x: bits_out=15'b110101111111101;
        15'b10x10x11111110x: bits_out=15'b101101111111101;
        15'b0x110x11111110x: bits_out=15'b011101111111101;
        15'b11110x11111110x: bits_out=15'b111101111111101;
        15'b10x0x111111110x: bits_out=15'b101011111111101;
        15'b0x10x111111110x: bits_out=15'b011011111111101;
        15'b1110x111111110x: bits_out=15'b111011111111101;
        15'b0x0x1111111110x: bits_out=15'b010111111111101;
        15'b110x1111111110x: bits_out=15'b110111111111101;
        15'b10x11111111110x: bits_out=15'b101111111111101;
        15'b0x111111111110x: bits_out=15'b011111111111101;
        15'b11111111111110x: bits_out=15'b111111111111101;
        15'b10x0x0x0x0x0x10: bits_out=15'b101010101010110;
        15'b0x10x0x0x0x0x10: bits_out=15'b011010101010110;
        15'b1110x0x0x0x0x10: bits_out=15'b111010101010110;
        15'b0x0x10x0x0x0x10: bits_out=15'b010110101010110;
        15'b110x10x0x0x0x10: bits_out=15'b110110101010110;
        15'b10x110x0x0x0x10: bits_out=15'b101110101010110;
        15'b0x1110x0x0x0x10: bits_out=15'b011110101010110;
        15'b111110x0x0x0x10: bits_out=15'b111110101010110;
        15'b0x0x0x10x0x0x10: bits_out=15'b010101101010110;
        15'b110x0x10x0x0x10: bits_out=15'b110101101010110;
        15'b10x10x10x0x0x10: bits_out=15'b101101101010110;
        15'b0x110x10x0x0x10: bits_out=15'b011101101010110;
        15'b11110x10x0x0x10: bits_out=15'b111101101010110;
        15'b10x0x110x0x0x10: bits_out=15'b101011101010110;
        15'b0x10x110x0x0x10: bits_out=15'b011011101010110;
        15'b1110x110x0x0x10: bits_out=15'b111011101010110;
        15'b0x0x1110x0x0x10: bits_out=15'b010111101010110;
        15'b110x1110x0x0x10: bits_out=15'b110111101010110;
        15'b10x11110x0x0x10: bits_out=15'b101111101010110;
        15'b0x111110x0x0x10: bits_out=15'b011111101010110;
        15'b11111110x0x0x10: bits_out=15'b111111101010110;
        15'b0x0x0x0x10x0x10: bits_out=15'b010101011010110;
        15'b110x0x0x10x0x10: bits_out=15'b110101011010110;
        15'b10x10x0x10x0x10: bits_out=15'b101101011010110;
        15'b0x110x0x10x0x10: bits_out=15'b011101011010110;
        15'b11110x0x10x0x10: bits_out=15'b111101011010110;
        15'b10x0x10x10x0x10: bits_out=15'b101011011010110;
        15'b0x10x10x10x0x10: bits_out=15'b011011011010110;
        15'b1110x10x10x0x10: bits_out=15'b111011011010110;
        15'b0x0x110x10x0x10: bits_out=15'b010111011010110;
        15'b110x110x10x0x10: bits_out=15'b110111011010110;
        15'b10x1110x10x0x10: bits_out=15'b101111011010110;
        15'b0x11110x10x0x10: bits_out=15'b011111011010110;
        15'b1111110x10x0x10: bits_out=15'b111111011010110;
        15'b10x0x0x110x0x10: bits_out=15'b101010111010110;
        15'b0x10x0x110x0x10: bits_out=15'b011010111010110;
        15'b1110x0x110x0x10: bits_out=15'b111010111010110;
        15'b0x0x10x110x0x10: bits_out=15'b010110111010110;
        15'b110x10x110x0x10: bits_out=15'b110110111010110;
        15'b10x110x110x0x10: bits_out=15'b101110111010110;
        15'b0x1110x110x0x10: bits_out=15'b011110111010110;
        15'b111110x110x0x10: bits_out=15'b111110111010110;
        15'b0x0x0x1110x0x10: bits_out=15'b010101111010110;
        15'b110x0x1110x0x10: bits_out=15'b110101111010110;
        15'b10x10x1110x0x10: bits_out=15'b101101111010110;
        15'b0x110x1110x0x10: bits_out=15'b011101111010110;
        15'b11110x1110x0x10: bits_out=15'b111101111010110;
        15'b10x0x11110x0x10: bits_out=15'b101011111010110;
        15'b0x10x11110x0x10: bits_out=15'b011011111010110;
        15'b1110x11110x0x10: bits_out=15'b111011111010110;
        15'b0x0x111110x0x10: bits_out=15'b010111111010110;
        15'b110x111110x0x10: bits_out=15'b110111111010110;
        15'b10x1111110x0x10: bits_out=15'b101111111010110;
        15'b0x11111110x0x10: bits_out=15'b011111111010110;
        15'b1111111110x0x10: bits_out=15'b111111111010110;
        15'b0x0x0x0x0x10x10: bits_out=15'b010101010110110;
        15'b110x0x0x0x10x10: bits_out=15'b110101010110110;
        15'b10x10x0x0x10x10: bits_out=15'b101101010110110;
        15'b0x110x0x0x10x10: bits_out=15'b011101010110110;
        15'b11110x0x0x10x10: bits_out=15'b111101010110110;
        15'b10x0x10x0x10x10: bits_out=15'b101011010110110;
        15'b0x10x10x0x10x10: bits_out=15'b011011010110110;
        15'b1110x10x0x10x10: bits_out=15'b111011010110110;
        15'b0x0x110x0x10x10: bits_out=15'b010111010110110;
        15'b110x110x0x10x10: bits_out=15'b110111010110110;
        15'b10x1110x0x10x10: bits_out=15'b101111010110110;
        15'b0x11110x0x10x10: bits_out=15'b011111010110110;
        15'b1111110x0x10x10: bits_out=15'b111111010110110;
        15'b10x0x0x10x10x10: bits_out=15'b101010110110110;
        15'b0x10x0x10x10x10: bits_out=15'b011010110110110;
        15'b1110x0x10x10x10: bits_out=15'b111010110110110;
        15'b0x0x10x10x10x10: bits_out=15'b010110110110110;
        15'b110x10x10x10x10: bits_out=15'b110110110110110;
        15'b10x110x10x10x10: bits_out=15'b101110110110110;
        15'b0x1110x10x10x10: bits_out=15'b011110110110110;
        15'b111110x10x10x10: bits_out=15'b111110110110110;
        15'b0x0x0x110x10x10: bits_out=15'b010101110110110;
        15'b110x0x110x10x10: bits_out=15'b110101110110110;
        15'b10x10x110x10x10: bits_out=15'b101101110110110;
        15'b0x110x110x10x10: bits_out=15'b011101110110110;
        15'b11110x110x10x10: bits_out=15'b111101110110110;
        15'b10x0x1110x10x10: bits_out=15'b101011110110110;
        15'b0x10x1110x10x10: bits_out=15'b011011110110110;
        15'b1110x1110x10x10: bits_out=15'b111011110110110;
        15'b0x0x11110x10x10: bits_out=15'b010111110110110;
        15'b110x11110x10x10: bits_out=15'b110111110110110;
        15'b10x111110x10x10: bits_out=15'b101111110110110;
        15'b0x1111110x10x10: bits_out=15'b011111110110110;
        15'b111111110x10x10: bits_out=15'b111111110110110;
        15'b10x0x0x0x110x10: bits_out=15'b101010101110110;
        15'b0x10x0x0x110x10: bits_out=15'b011010101110110;
        15'b1110x0x0x110x10: bits_out=15'b111010101110110;
        15'b0x0x10x0x110x10: bits_out=15'b010110101110110;
        15'b110x10x0x110x10: bits_out=15'b110110101110110;
        15'b10x110x0x110x10: bits_out=15'b101110101110110;
        15'b0x1110x0x110x10: bits_out=15'b011110101110110;
        15'b111110x0x110x10: bits_out=15'b111110101110110;
        15'b0x0x0x10x110x10: bits_out=15'b010101101110110;
        15'b110x0x10x110x10: bits_out=15'b110101101110110;
        15'b10x10x10x110x10: bits_out=15'b101101101110110;
        15'b0x110x10x110x10: bits_out=15'b011101101110110;
        15'b11110x10x110x10: bits_out=15'b111101101110110;
        15'b10x0x110x110x10: bits_out=15'b101011101110110;
        15'b0x10x110x110x10: bits_out=15'b011011101110110;
        15'b1110x110x110x10: bits_out=15'b111011101110110;
        15'b0x0x1110x110x10: bits_out=15'b010111101110110;
        15'b110x1110x110x10: bits_out=15'b110111101110110;
        15'b10x11110x110x10: bits_out=15'b101111101110110;
        15'b0x111110x110x10: bits_out=15'b011111101110110;
        15'b11111110x110x10: bits_out=15'b111111101110110;
        15'b0x0x0x0x1110x10: bits_out=15'b010101011110110;
        15'b110x0x0x1110x10: bits_out=15'b110101011110110;
        15'b10x10x0x1110x10: bits_out=15'b101101011110110;
        15'b0x110x0x1110x10: bits_out=15'b011101011110110;
        15'b11110x0x1110x10: bits_out=15'b111101011110110;
        15'b10x0x10x1110x10: bits_out=15'b101011011110110;
        15'b0x10x10x1110x10: bits_out=15'b011011011110110;
        15'b1110x10x1110x10: bits_out=15'b111011011110110;
        15'b0x0x110x1110x10: bits_out=15'b010111011110110;
        15'b110x110x1110x10: bits_out=15'b110111011110110;
        15'b10x1110x1110x10: bits_out=15'b101111011110110;
        15'b0x11110x1110x10: bits_out=15'b011111011110110;
        15'b1111110x1110x10: bits_out=15'b111111011110110;
        15'b10x0x0x11110x10: bits_out=15'b101010111110110;
        15'b0x10x0x11110x10: bits_out=15'b011010111110110;
        15'b1110x0x11110x10: bits_out=15'b111010111110110;
        15'b0x0x10x11110x10: bits_out=15'b010110111110110;
        15'b110x10x11110x10: bits_out=15'b110110111110110;
        15'b10x110x11110x10: bits_out=15'b101110111110110;
        15'b0x1110x11110x10: bits_out=15'b011110111110110;
        15'b111110x11110x10: bits_out=15'b111110111110110;
        15'b0x0x0x111110x10: bits_out=15'b010101111110110;
        15'b110x0x111110x10: bits_out=15'b110101111110110;
        15'b10x10x111110x10: bits_out=15'b101101111110110;
        15'b0x110x111110x10: bits_out=15'b011101111110110;
        15'b11110x111110x10: bits_out=15'b111101111110110;
        15'b10x0x1111110x10: bits_out=15'b101011111110110;
        15'b0x10x1111110x10: bits_out=15'b011011111110110;
        15'b1110x1111110x10: bits_out=15'b111011111110110;
        15'b0x0x11111110x10: bits_out=15'b010111111110110;
        15'b110x11111110x10: bits_out=15'b110111111110110;
        15'b10x111111110x10: bits_out=15'b101111111110110;
        15'b0x1111111110x10: bits_out=15'b011111111110110;
        15'b111111111110x10: bits_out=15'b111111111110110;
        15'b0x0x0x0x0x0x110: bits_out=15'b010101010101110;
        15'b110x0x0x0x0x110: bits_out=15'b110101010101110;
        15'b10x10x0x0x0x110: bits_out=15'b101101010101110;
        15'b0x110x0x0x0x110: bits_out=15'b011101010101110;
        15'b11110x0x0x0x110: bits_out=15'b111101010101110;
        15'b10x0x10x0x0x110: bits_out=15'b101011010101110;
        15'b0x10x10x0x0x110: bits_out=15'b011011010101110;
        15'b1110x10x0x0x110: bits_out=15'b111011010101110;
        15'b0x0x110x0x0x110: bits_out=15'b010111010101110;
        15'b110x110x0x0x110: bits_out=15'b110111010101110;
        15'b10x1110x0x0x110: bits_out=15'b101111010101110;
        15'b0x11110x0x0x110: bits_out=15'b011111010101110;
        15'b1111110x0x0x110: bits_out=15'b111111010101110;
        15'b10x0x0x10x0x110: bits_out=15'b101010110101110;
        15'b0x10x0x10x0x110: bits_out=15'b011010110101110;
        15'b1110x0x10x0x110: bits_out=15'b111010110101110;
        15'b0x0x10x10x0x110: bits_out=15'b010110110101110;
        15'b110x10x10x0x110: bits_out=15'b110110110101110;
        15'b10x110x10x0x110: bits_out=15'b101110110101110;
        15'b0x1110x10x0x110: bits_out=15'b011110110101110;
        15'b111110x10x0x110: bits_out=15'b111110110101110;
        15'b0x0x0x110x0x110: bits_out=15'b010101110101110;
        15'b110x0x110x0x110: bits_out=15'b110101110101110;
        15'b10x10x110x0x110: bits_out=15'b101101110101110;
        15'b0x110x110x0x110: bits_out=15'b011101110101110;
        15'b11110x110x0x110: bits_out=15'b111101110101110;
        15'b10x0x1110x0x110: bits_out=15'b101011110101110;
        15'b0x10x1110x0x110: bits_out=15'b011011110101110;
        15'b1110x1110x0x110: bits_out=15'b111011110101110;
        15'b0x0x11110x0x110: bits_out=15'b010111110101110;
        15'b110x11110x0x110: bits_out=15'b110111110101110;
        15'b10x111110x0x110: bits_out=15'b101111110101110;
        15'b0x1111110x0x110: bits_out=15'b011111110101110;
        15'b111111110x0x110: bits_out=15'b111111110101110;
        15'b10x0x0x0x10x110: bits_out=15'b101010101101110;
        15'b0x10x0x0x10x110: bits_out=15'b011010101101110;
        15'b1110x0x0x10x110: bits_out=15'b111010101101110;
        15'b0x0x10x0x10x110: bits_out=15'b010110101101110;
        15'b110x10x0x10x110: bits_out=15'b110110101101110;
        15'b10x110x0x10x110: bits_out=15'b101110101101110;
        15'b0x1110x0x10x110: bits_out=15'b011110101101110;
        15'b111110x0x10x110: bits_out=15'b111110101101110;
        15'b0x0x0x10x10x110: bits_out=15'b010101101101110;
        15'b110x0x10x10x110: bits_out=15'b110101101101110;
        15'b10x10x10x10x110: bits_out=15'b101101101101110;
        15'b0x110x10x10x110: bits_out=15'b011101101101110;
        15'b11110x10x10x110: bits_out=15'b111101101101110;
        15'b10x0x110x10x110: bits_out=15'b101011101101110;
        15'b0x10x110x10x110: bits_out=15'b011011101101110;
        15'b1110x110x10x110: bits_out=15'b111011101101110;
        15'b0x0x1110x10x110: bits_out=15'b010111101101110;
        15'b110x1110x10x110: bits_out=15'b110111101101110;
        15'b10x11110x10x110: bits_out=15'b101111101101110;
        15'b0x111110x10x110: bits_out=15'b011111101101110;
        15'b11111110x10x110: bits_out=15'b111111101101110;
        15'b0x0x0x0x110x110: bits_out=15'b010101011101110;
        15'b110x0x0x110x110: bits_out=15'b110101011101110;
        15'b10x10x0x110x110: bits_out=15'b101101011101110;
        15'b0x110x0x110x110: bits_out=15'b011101011101110;
        15'b11110x0x110x110: bits_out=15'b111101011101110;
        15'b10x0x10x110x110: bits_out=15'b101011011101110;
        15'b0x10x10x110x110: bits_out=15'b011011011101110;
        15'b1110x10x110x110: bits_out=15'b111011011101110;
        15'b0x0x110x110x110: bits_out=15'b010111011101110;
        15'b110x110x110x110: bits_out=15'b110111011101110;
        15'b10x1110x110x110: bits_out=15'b101111011101110;
        15'b0x11110x110x110: bits_out=15'b011111011101110;
        15'b1111110x110x110: bits_out=15'b111111011101110;
        15'b10x0x0x1110x110: bits_out=15'b101010111101110;
        15'b0x10x0x1110x110: bits_out=15'b011010111101110;
        15'b1110x0x1110x110: bits_out=15'b111010111101110;
        15'b0x0x10x1110x110: bits_out=15'b010110111101110;
        15'b110x10x1110x110: bits_out=15'b110110111101110;
        15'b10x110x1110x110: bits_out=15'b101110111101110;
        15'b0x1110x1110x110: bits_out=15'b011110111101110;
        15'b111110x1110x110: bits_out=15'b111110111101110;
        15'b0x0x0x11110x110: bits_out=15'b010101111101110;
        15'b110x0x11110x110: bits_out=15'b110101111101110;
        15'b10x10x11110x110: bits_out=15'b101101111101110;
        15'b0x110x11110x110: bits_out=15'b011101111101110;
        15'b11110x11110x110: bits_out=15'b111101111101110;
        15'b10x0x111110x110: bits_out=15'b101011111101110;
        15'b0x10x111110x110: bits_out=15'b011011111101110;
        15'b1110x111110x110: bits_out=15'b111011111101110;
        15'b0x0x1111110x110: bits_out=15'b010111111101110;
        15'b110x1111110x110: bits_out=15'b110111111101110;
        15'b10x11111110x110: bits_out=15'b101111111101110;
        15'b0x111111110x110: bits_out=15'b011111111101110;
        15'b11111111110x110: bits_out=15'b111111111101110;
        15'b10x0x0x0x0x1110: bits_out=15'b101010101011110;
        15'b0x10x0x0x0x1110: bits_out=15'b011010101011110;
        15'b1110x0x0x0x1110: bits_out=15'b111010101011110;
        15'b0x0x10x0x0x1110: bits_out=15'b010110101011110;
        15'b110x10x0x0x1110: bits_out=15'b110110101011110;
        15'b10x110x0x0x1110: bits_out=15'b101110101011110;
        15'b0x1110x0x0x1110: bits_out=15'b011110101011110;
        15'b111110x0x0x1110: bits_out=15'b111110101011110;
        15'b0x0x0x10x0x1110: bits_out=15'b010101101011110;
        15'b110x0x10x0x1110: bits_out=15'b110101101011110;
        15'b10x10x10x0x1110: bits_out=15'b101101101011110;
        15'b0x110x10x0x1110: bits_out=15'b011101101011110;
        15'b11110x10x0x1110: bits_out=15'b111101101011110;
        15'b10x0x110x0x1110: bits_out=15'b101011101011110;
        15'b0x10x110x0x1110: bits_out=15'b011011101011110;
        15'b1110x110x0x1110: bits_out=15'b111011101011110;
        15'b0x0x1110x0x1110: bits_out=15'b010111101011110;
        15'b110x1110x0x1110: bits_out=15'b110111101011110;
        15'b10x11110x0x1110: bits_out=15'b101111101011110;
        15'b0x111110x0x1110: bits_out=15'b011111101011110;
        15'b11111110x0x1110: bits_out=15'b111111101011110;
        15'b0x0x0x0x10x1110: bits_out=15'b010101011011110;
        15'b110x0x0x10x1110: bits_out=15'b110101011011110;
        15'b10x10x0x10x1110: bits_out=15'b101101011011110;
        15'b0x110x0x10x1110: bits_out=15'b011101011011110;
        15'b11110x0x10x1110: bits_out=15'b111101011011110;
        15'b10x0x10x10x1110: bits_out=15'b101011011011110;
        15'b0x10x10x10x1110: bits_out=15'b011011011011110;
        15'b1110x10x10x1110: bits_out=15'b111011011011110;
        15'b0x0x110x10x1110: bits_out=15'b010111011011110;
        15'b110x110x10x1110: bits_out=15'b110111011011110;
        15'b10x1110x10x1110: bits_out=15'b101111011011110;
        15'b0x11110x10x1110: bits_out=15'b011111011011110;
        15'b1111110x10x1110: bits_out=15'b111111011011110;
        15'b10x0x0x110x1110: bits_out=15'b101010111011110;
        15'b0x10x0x110x1110: bits_out=15'b011010111011110;
        15'b1110x0x110x1110: bits_out=15'b111010111011110;
        15'b0x0x10x110x1110: bits_out=15'b010110111011110;
        15'b110x10x110x1110: bits_out=15'b110110111011110;
        15'b10x110x110x1110: bits_out=15'b101110111011110;
        15'b0x1110x110x1110: bits_out=15'b011110111011110;
        15'b111110x110x1110: bits_out=15'b111110111011110;
        15'b0x0x0x1110x1110: bits_out=15'b010101111011110;
        15'b110x0x1110x1110: bits_out=15'b110101111011110;
        15'b10x10x1110x1110: bits_out=15'b101101111011110;
        15'b0x110x1110x1110: bits_out=15'b011101111011110;
        15'b11110x1110x1110: bits_out=15'b111101111011110;
        15'b10x0x11110x1110: bits_out=15'b101011111011110;
        15'b0x10x11110x1110: bits_out=15'b011011111011110;
        15'b1110x11110x1110: bits_out=15'b111011111011110;
        15'b0x0x111110x1110: bits_out=15'b010111111011110;
        15'b110x111110x1110: bits_out=15'b110111111011110;
        15'b10x1111110x1110: bits_out=15'b101111111011110;
        15'b0x11111110x1110: bits_out=15'b011111111011110;
        15'b1111111110x1110: bits_out=15'b111111111011110;
        15'b0x0x0x0x0x11110: bits_out=15'b010101010111110;
        15'b110x0x0x0x11110: bits_out=15'b110101010111110;
        15'b10x10x0x0x11110: bits_out=15'b101101010111110;
        15'b0x110x0x0x11110: bits_out=15'b011101010111110;
        15'b11110x0x0x11110: bits_out=15'b111101010111110;
        15'b10x0x10x0x11110: bits_out=15'b101011010111110;
        15'b0x10x10x0x11110: bits_out=15'b011011010111110;
        15'b1110x10x0x11110: bits_out=15'b111011010111110;
        15'b0x0x110x0x11110: bits_out=15'b010111010111110;
        15'b110x110x0x11110: bits_out=15'b110111010111110;
        15'b10x1110x0x11110: bits_out=15'b101111010111110;
        15'b0x11110x0x11110: bits_out=15'b011111010111110;
        15'b1111110x0x11110: bits_out=15'b111111010111110;
        15'b10x0x0x10x11110: bits_out=15'b101010110111110;
        15'b0x10x0x10x11110: bits_out=15'b011010110111110;
        15'b1110x0x10x11110: bits_out=15'b111010110111110;
        15'b0x0x10x10x11110: bits_out=15'b010110110111110;
        15'b110x10x10x11110: bits_out=15'b110110110111110;
        15'b10x110x10x11110: bits_out=15'b101110110111110;
        15'b0x1110x10x11110: bits_out=15'b011110110111110;
        15'b111110x10x11110: bits_out=15'b111110110111110;
        15'b0x0x0x110x11110: bits_out=15'b010101110111110;
        15'b110x0x110x11110: bits_out=15'b110101110111110;
        15'b10x10x110x11110: bits_out=15'b101101110111110;
        15'b0x110x110x11110: bits_out=15'b011101110111110;
        15'b11110x110x11110: bits_out=15'b111101110111110;
        15'b10x0x1110x11110: bits_out=15'b101011110111110;
        15'b0x10x1110x11110: bits_out=15'b011011110111110;
        15'b1110x1110x11110: bits_out=15'b111011110111110;
        15'b0x0x11110x11110: bits_out=15'b010111110111110;
        15'b110x11110x11110: bits_out=15'b110111110111110;
        15'b10x111110x11110: bits_out=15'b101111110111110;
        15'b0x1111110x11110: bits_out=15'b011111110111110;
        15'b111111110x11110: bits_out=15'b111111110111110;
        15'b10x0x0x0x111110: bits_out=15'b101010101111110;
        15'b0x10x0x0x111110: bits_out=15'b011010101111110;
        15'b1110x0x0x111110: bits_out=15'b111010101111110;
        15'b0x0x10x0x111110: bits_out=15'b010110101111110;
        15'b110x10x0x111110: bits_out=15'b110110101111110;
        15'b10x110x0x111110: bits_out=15'b101110101111110;
        15'b0x1110x0x111110: bits_out=15'b011110101111110;
        15'b111110x0x111110: bits_out=15'b111110101111110;
        15'b0x0x0x10x111110: bits_out=15'b010101101111110;
        15'b110x0x10x111110: bits_out=15'b110101101111110;
        15'b10x10x10x111110: bits_out=15'b101101101111110;
        15'b0x110x10x111110: bits_out=15'b011101101111110;
        15'b11110x10x111110: bits_out=15'b111101101111110;
        15'b10x0x110x111110: bits_out=15'b101011101111110;
        15'b0x10x110x111110: bits_out=15'b011011101111110;
        15'b1110x110x111110: bits_out=15'b111011101111110;
        15'b0x0x1110x111110: bits_out=15'b010111101111110;
        15'b110x1110x111110: bits_out=15'b110111101111110;
        15'b10x11110x111110: bits_out=15'b101111101111110;
        15'b0x111110x111110: bits_out=15'b011111101111110;
        15'b11111110x111110: bits_out=15'b111111101111110;
        15'b0x0x0x0x1111110: bits_out=15'b010101011111110;
        15'b110x0x0x1111110: bits_out=15'b110101011111110;
        15'b10x10x0x1111110: bits_out=15'b101101011111110;
        15'b0x110x0x1111110: bits_out=15'b011101011111110;
        15'b11110x0x1111110: bits_out=15'b111101011111110;
        15'b10x0x10x1111110: bits_out=15'b101011011111110;
        15'b0x10x10x1111110: bits_out=15'b011011011111110;
        15'b1110x10x1111110: bits_out=15'b111011011111110;
        15'b0x0x110x1111110: bits_out=15'b010111011111110;
        15'b110x110x1111110: bits_out=15'b110111011111110;
        15'b10x1110x1111110: bits_out=15'b101111011111110;
        15'b0x11110x1111110: bits_out=15'b011111011111110;
        15'b1111110x1111110: bits_out=15'b111111011111110;
        15'b10x0x0x11111110: bits_out=15'b101010111111110;
        15'b0x10x0x11111110: bits_out=15'b011010111111110;
        15'b1110x0x11111110: bits_out=15'b111010111111110;
        15'b0x0x10x11111110: bits_out=15'b010110111111110;
        15'b110x10x11111110: bits_out=15'b110110111111110;
        15'b10x110x11111110: bits_out=15'b101110111111110;
        15'b0x1110x11111110: bits_out=15'b011110111111110;
        15'b111110x11111110: bits_out=15'b111110111111110;
        15'b0x0x0x111111110: bits_out=15'b010101111111110;
        15'b110x0x111111110: bits_out=15'b110101111111110;
        15'b10x10x111111110: bits_out=15'b101101111111110;
        15'b0x110x111111110: bits_out=15'b011101111111110;
        15'b11110x111111110: bits_out=15'b111101111111110;
        15'b10x0x1111111110: bits_out=15'b101011111111110;
        15'b0x10x1111111110: bits_out=15'b011011111111110;
        15'b1110x1111111110: bits_out=15'b111011111111110;
        15'b0x0x11111111110: bits_out=15'b010111111111110;
        15'b110x11111111110: bits_out=15'b110111111111110;
        15'b10x111111111110: bits_out=15'b101111111111110;
        15'b0x1111111111110: bits_out=15'b011111111111110;
        15'b111111111111110: bits_out=15'b111111111111110;
        15'b0x0x0x0x0x0x0x1: bits_out=15'b010101010101011;
        15'b110x0x0x0x0x0x1: bits_out=15'b110101010101011;
        15'b10x10x0x0x0x0x1: bits_out=15'b101101010101011;
        15'b0x110x0x0x0x0x1: bits_out=15'b011101010101011;
        15'b11110x0x0x0x0x1: bits_out=15'b111101010101011;
        15'b10x0x10x0x0x0x1: bits_out=15'b101011010101011;
        15'b0x10x10x0x0x0x1: bits_out=15'b011011010101011;
        15'b1110x10x0x0x0x1: bits_out=15'b111011010101011;
        15'b0x0x110x0x0x0x1: bits_out=15'b010111010101011;
        15'b110x110x0x0x0x1: bits_out=15'b110111010101011;
        15'b10x1110x0x0x0x1: bits_out=15'b101111010101011;
        15'b0x11110x0x0x0x1: bits_out=15'b011111010101011;
        15'b1111110x0x0x0x1: bits_out=15'b111111010101011;
        15'b10x0x0x10x0x0x1: bits_out=15'b101010110101011;
        15'b0x10x0x10x0x0x1: bits_out=15'b011010110101011;
        15'b1110x0x10x0x0x1: bits_out=15'b111010110101011;
        15'b0x0x10x10x0x0x1: bits_out=15'b010110110101011;
        15'b110x10x10x0x0x1: bits_out=15'b110110110101011;
        15'b10x110x10x0x0x1: bits_out=15'b101110110101011;
        15'b0x1110x10x0x0x1: bits_out=15'b011110110101011;
        15'b111110x10x0x0x1: bits_out=15'b111110110101011;
        15'b0x0x0x110x0x0x1: bits_out=15'b010101110101011;
        15'b110x0x110x0x0x1: bits_out=15'b110101110101011;
        15'b10x10x110x0x0x1: bits_out=15'b101101110101011;
        15'b0x110x110x0x0x1: bits_out=15'b011101110101011;
        15'b11110x110x0x0x1: bits_out=15'b111101110101011;
        15'b10x0x1110x0x0x1: bits_out=15'b101011110101011;
        15'b0x10x1110x0x0x1: bits_out=15'b011011110101011;
        15'b1110x1110x0x0x1: bits_out=15'b111011110101011;
        15'b0x0x11110x0x0x1: bits_out=15'b010111110101011;
        15'b110x11110x0x0x1: bits_out=15'b110111110101011;
        15'b10x111110x0x0x1: bits_out=15'b101111110101011;
        15'b0x1111110x0x0x1: bits_out=15'b011111110101011;
        15'b111111110x0x0x1: bits_out=15'b111111110101011;
        15'b10x0x0x0x10x0x1: bits_out=15'b101010101101011;
        15'b0x10x0x0x10x0x1: bits_out=15'b011010101101011;
        15'b1110x0x0x10x0x1: bits_out=15'b111010101101011;
        15'b0x0x10x0x10x0x1: bits_out=15'b010110101101011;
        15'b110x10x0x10x0x1: bits_out=15'b110110101101011;
        15'b10x110x0x10x0x1: bits_out=15'b101110101101011;
        15'b0x1110x0x10x0x1: bits_out=15'b011110101101011;
        15'b111110x0x10x0x1: bits_out=15'b111110101101011;
        15'b0x0x0x10x10x0x1: bits_out=15'b010101101101011;
        15'b110x0x10x10x0x1: bits_out=15'b110101101101011;
        15'b10x10x10x10x0x1: bits_out=15'b101101101101011;
        15'b0x110x10x10x0x1: bits_out=15'b011101101101011;
        15'b11110x10x10x0x1: bits_out=15'b111101101101011;
        15'b10x0x110x10x0x1: bits_out=15'b101011101101011;
        15'b0x10x110x10x0x1: bits_out=15'b011011101101011;
        15'b1110x110x10x0x1: bits_out=15'b111011101101011;
        15'b0x0x1110x10x0x1: bits_out=15'b010111101101011;
        15'b110x1110x10x0x1: bits_out=15'b110111101101011;
        15'b10x11110x10x0x1: bits_out=15'b101111101101011;
        15'b0x111110x10x0x1: bits_out=15'b011111101101011;
        15'b11111110x10x0x1: bits_out=15'b111111101101011;
        15'b0x0x0x0x110x0x1: bits_out=15'b010101011101011;
        15'b110x0x0x110x0x1: bits_out=15'b110101011101011;
        15'b10x10x0x110x0x1: bits_out=15'b101101011101011;
        15'b0x110x0x110x0x1: bits_out=15'b011101011101011;
        15'b11110x0x110x0x1: bits_out=15'b111101011101011;
        15'b10x0x10x110x0x1: bits_out=15'b101011011101011;
        15'b0x10x10x110x0x1: bits_out=15'b011011011101011;
        15'b1110x10x110x0x1: bits_out=15'b111011011101011;
        15'b0x0x110x110x0x1: bits_out=15'b010111011101011;
        15'b110x110x110x0x1: bits_out=15'b110111011101011;
        15'b10x1110x110x0x1: bits_out=15'b101111011101011;
        15'b0x11110x110x0x1: bits_out=15'b011111011101011;
        15'b1111110x110x0x1: bits_out=15'b111111011101011;
        15'b10x0x0x1110x0x1: bits_out=15'b101010111101011;
        15'b0x10x0x1110x0x1: bits_out=15'b011010111101011;
        15'b1110x0x1110x0x1: bits_out=15'b111010111101011;
        15'b0x0x10x1110x0x1: bits_out=15'b010110111101011;
        15'b110x10x1110x0x1: bits_out=15'b110110111101011;
        15'b10x110x1110x0x1: bits_out=15'b101110111101011;
        15'b0x1110x1110x0x1: bits_out=15'b011110111101011;
        15'b111110x1110x0x1: bits_out=15'b111110111101011;
        15'b0x0x0x11110x0x1: bits_out=15'b010101111101011;
        15'b110x0x11110x0x1: bits_out=15'b110101111101011;
        15'b10x10x11110x0x1: bits_out=15'b101101111101011;
        15'b0x110x11110x0x1: bits_out=15'b011101111101011;
        15'b11110x11110x0x1: bits_out=15'b111101111101011;
        15'b10x0x111110x0x1: bits_out=15'b101011111101011;
        15'b0x10x111110x0x1: bits_out=15'b011011111101011;
        15'b1110x111110x0x1: bits_out=15'b111011111101011;
        15'b0x0x1111110x0x1: bits_out=15'b010111111101011;
        15'b110x1111110x0x1: bits_out=15'b110111111101011;
        15'b10x11111110x0x1: bits_out=15'b101111111101011;
        15'b0x111111110x0x1: bits_out=15'b011111111101011;
        15'b11111111110x0x1: bits_out=15'b111111111101011;
        15'b10x0x0x0x0x10x1: bits_out=15'b101010101011011;
        15'b0x10x0x0x0x10x1: bits_out=15'b011010101011011;
        15'b1110x0x0x0x10x1: bits_out=15'b111010101011011;
        15'b0x0x10x0x0x10x1: bits_out=15'b010110101011011;
        15'b110x10x0x0x10x1: bits_out=15'b110110101011011;
        15'b10x110x0x0x10x1: bits_out=15'b101110101011011;
        15'b0x1110x0x0x10x1: bits_out=15'b011110101011011;
        15'b111110x0x0x10x1: bits_out=15'b111110101011011;
        15'b0x0x0x10x0x10x1: bits_out=15'b010101101011011;
        15'b110x0x10x0x10x1: bits_out=15'b110101101011011;
        15'b10x10x10x0x10x1: bits_out=15'b101101101011011;
        15'b0x110x10x0x10x1: bits_out=15'b011101101011011;
        15'b11110x10x0x10x1: bits_out=15'b111101101011011;
        15'b10x0x110x0x10x1: bits_out=15'b101011101011011;
        15'b0x10x110x0x10x1: bits_out=15'b011011101011011;
        15'b1110x110x0x10x1: bits_out=15'b111011101011011;
        15'b0x0x1110x0x10x1: bits_out=15'b010111101011011;
        15'b110x1110x0x10x1: bits_out=15'b110111101011011;
        15'b10x11110x0x10x1: bits_out=15'b101111101011011;
        15'b0x111110x0x10x1: bits_out=15'b011111101011011;
        15'b11111110x0x10x1: bits_out=15'b111111101011011;
        15'b0x0x0x0x10x10x1: bits_out=15'b010101011011011;
        15'b110x0x0x10x10x1: bits_out=15'b110101011011011;
        15'b10x10x0x10x10x1: bits_out=15'b101101011011011;
        15'b0x110x0x10x10x1: bits_out=15'b011101011011011;
        15'b11110x0x10x10x1: bits_out=15'b111101011011011;
        15'b10x0x10x10x10x1: bits_out=15'b101011011011011;
        15'b0x10x10x10x10x1: bits_out=15'b011011011011011;
        15'b1110x10x10x10x1: bits_out=15'b111011011011011;
        15'b0x0x110x10x10x1: bits_out=15'b010111011011011;
        15'b110x110x10x10x1: bits_out=15'b110111011011011;
        15'b10x1110x10x10x1: bits_out=15'b101111011011011;
        15'b0x11110x10x10x1: bits_out=15'b011111011011011;
        15'b1111110x10x10x1: bits_out=15'b111111011011011;
        15'b10x0x0x110x10x1: bits_out=15'b101010111011011;
        15'b0x10x0x110x10x1: bits_out=15'b011010111011011;
        15'b1110x0x110x10x1: bits_out=15'b111010111011011;
        15'b0x0x10x110x10x1: bits_out=15'b010110111011011;
        15'b110x10x110x10x1: bits_out=15'b110110111011011;
        15'b10x110x110x10x1: bits_out=15'b101110111011011;
        15'b0x1110x110x10x1: bits_out=15'b011110111011011;
        15'b111110x110x10x1: bits_out=15'b111110111011011;
        15'b0x0x0x1110x10x1: bits_out=15'b010101111011011;
        15'b110x0x1110x10x1: bits_out=15'b110101111011011;
        15'b10x10x1110x10x1: bits_out=15'b101101111011011;
        15'b0x110x1110x10x1: bits_out=15'b011101111011011;
        15'b11110x1110x10x1: bits_out=15'b111101111011011;
        15'b10x0x11110x10x1: bits_out=15'b101011111011011;
        15'b0x10x11110x10x1: bits_out=15'b011011111011011;
        15'b1110x11110x10x1: bits_out=15'b111011111011011;
        15'b0x0x111110x10x1: bits_out=15'b010111111011011;
        15'b110x111110x10x1: bits_out=15'b110111111011011;
        15'b10x1111110x10x1: bits_out=15'b101111111011011;
        15'b0x11111110x10x1: bits_out=15'b011111111011011;
        15'b1111111110x10x1: bits_out=15'b111111111011011;
        15'b0x0x0x0x0x110x1: bits_out=15'b010101010111011;
        15'b110x0x0x0x110x1: bits_out=15'b110101010111011;
        15'b10x10x0x0x110x1: bits_out=15'b101101010111011;
        15'b0x110x0x0x110x1: bits_out=15'b011101010111011;
        15'b11110x0x0x110x1: bits_out=15'b111101010111011;
        15'b10x0x10x0x110x1: bits_out=15'b101011010111011;
        15'b0x10x10x0x110x1: bits_out=15'b011011010111011;
        15'b1110x10x0x110x1: bits_out=15'b111011010111011;
        15'b0x0x110x0x110x1: bits_out=15'b010111010111011;
        15'b110x110x0x110x1: bits_out=15'b110111010111011;
        15'b10x1110x0x110x1: bits_out=15'b101111010111011;
        15'b0x11110x0x110x1: bits_out=15'b011111010111011;
        15'b1111110x0x110x1: bits_out=15'b111111010111011;
        15'b10x0x0x10x110x1: bits_out=15'b101010110111011;
        15'b0x10x0x10x110x1: bits_out=15'b011010110111011;
        15'b1110x0x10x110x1: bits_out=15'b111010110111011;
        15'b0x0x10x10x110x1: bits_out=15'b010110110111011;
        15'b110x10x10x110x1: bits_out=15'b110110110111011;
        15'b10x110x10x110x1: bits_out=15'b101110110111011;
        15'b0x1110x10x110x1: bits_out=15'b011110110111011;
        15'b111110x10x110x1: bits_out=15'b111110110111011;
        15'b0x0x0x110x110x1: bits_out=15'b010101110111011;
        15'b110x0x110x110x1: bits_out=15'b110101110111011;
        15'b10x10x110x110x1: bits_out=15'b101101110111011;
        15'b0x110x110x110x1: bits_out=15'b011101110111011;
        15'b11110x110x110x1: bits_out=15'b111101110111011;
        15'b10x0x1110x110x1: bits_out=15'b101011110111011;
        15'b0x10x1110x110x1: bits_out=15'b011011110111011;
        15'b1110x1110x110x1: bits_out=15'b111011110111011;
        15'b0x0x11110x110x1: bits_out=15'b010111110111011;
        15'b110x11110x110x1: bits_out=15'b110111110111011;
        15'b10x111110x110x1: bits_out=15'b101111110111011;
        15'b0x1111110x110x1: bits_out=15'b011111110111011;
        15'b111111110x110x1: bits_out=15'b111111110111011;
        15'b10x0x0x0x1110x1: bits_out=15'b101010101111011;
        15'b0x10x0x0x1110x1: bits_out=15'b011010101111011;
        15'b1110x0x0x1110x1: bits_out=15'b111010101111011;
        15'b0x0x10x0x1110x1: bits_out=15'b010110101111011;
        15'b110x10x0x1110x1: bits_out=15'b110110101111011;
        15'b10x110x0x1110x1: bits_out=15'b101110101111011;
        15'b0x1110x0x1110x1: bits_out=15'b011110101111011;
        15'b111110x0x1110x1: bits_out=15'b111110101111011;
        15'b0x0x0x10x1110x1: bits_out=15'b010101101111011;
        15'b110x0x10x1110x1: bits_out=15'b110101101111011;
        15'b10x10x10x1110x1: bits_out=15'b101101101111011;
        15'b0x110x10x1110x1: bits_out=15'b011101101111011;
        15'b11110x10x1110x1: bits_out=15'b111101101111011;
        15'b10x0x110x1110x1: bits_out=15'b101011101111011;
        15'b0x10x110x1110x1: bits_out=15'b011011101111011;
        15'b1110x110x1110x1: bits_out=15'b111011101111011;
        15'b0x0x1110x1110x1: bits_out=15'b010111101111011;
        15'b110x1110x1110x1: bits_out=15'b110111101111011;
        15'b10x11110x1110x1: bits_out=15'b101111101111011;
        15'b0x111110x1110x1: bits_out=15'b011111101111011;
        15'b11111110x1110x1: bits_out=15'b111111101111011;
        15'b0x0x0x0x11110x1: bits_out=15'b010101011111011;
        15'b110x0x0x11110x1: bits_out=15'b110101011111011;
        15'b10x10x0x11110x1: bits_out=15'b101101011111011;
        15'b0x110x0x11110x1: bits_out=15'b011101011111011;
        15'b11110x0x11110x1: bits_out=15'b111101011111011;
        15'b10x0x10x11110x1: bits_out=15'b101011011111011;
        15'b0x10x10x11110x1: bits_out=15'b011011011111011;
        15'b1110x10x11110x1: bits_out=15'b111011011111011;
        15'b0x0x110x11110x1: bits_out=15'b010111011111011;
        15'b110x110x11110x1: bits_out=15'b110111011111011;
        15'b10x1110x11110x1: bits_out=15'b101111011111011;
        15'b0x11110x11110x1: bits_out=15'b011111011111011;
        15'b1111110x11110x1: bits_out=15'b111111011111011;
        15'b10x0x0x111110x1: bits_out=15'b101010111111011;
        15'b0x10x0x111110x1: bits_out=15'b011010111111011;
        15'b1110x0x111110x1: bits_out=15'b111010111111011;
        15'b0x0x10x111110x1: bits_out=15'b010110111111011;
        15'b110x10x111110x1: bits_out=15'b110110111111011;
        15'b10x110x111110x1: bits_out=15'b101110111111011;
        15'b0x1110x111110x1: bits_out=15'b011110111111011;
        15'b111110x111110x1: bits_out=15'b111110111111011;
        15'b0x0x0x1111110x1: bits_out=15'b010101111111011;
        15'b110x0x1111110x1: bits_out=15'b110101111111011;
        15'b10x10x1111110x1: bits_out=15'b101101111111011;
        15'b0x110x1111110x1: bits_out=15'b011101111111011;
        15'b11110x1111110x1: bits_out=15'b111101111111011;
        15'b10x0x11111110x1: bits_out=15'b101011111111011;
        15'b0x10x11111110x1: bits_out=15'b011011111111011;
        15'b1110x11111110x1: bits_out=15'b111011111111011;
        15'b0x0x111111110x1: bits_out=15'b010111111111011;
        15'b110x111111110x1: bits_out=15'b110111111111011;
        15'b10x1111111110x1: bits_out=15'b101111111111011;
        15'b0x11111111110x1: bits_out=15'b011111111111011;
        15'b1111111111110x1: bits_out=15'b111111111111011;
        15'b10x0x0x0x0x0x11: bits_out=15'b101010101010111;
        15'b0x10x0x0x0x0x11: bits_out=15'b011010101010111;
        15'b1110x0x0x0x0x11: bits_out=15'b111010101010111;
        15'b0x0x10x0x0x0x11: bits_out=15'b010110101010111;
        15'b110x10x0x0x0x11: bits_out=15'b110110101010111;
        15'b10x110x0x0x0x11: bits_out=15'b101110101010111;
        15'b0x1110x0x0x0x11: bits_out=15'b011110101010111;
        15'b111110x0x0x0x11: bits_out=15'b111110101010111;
        15'b0x0x0x10x0x0x11: bits_out=15'b010101101010111;
        15'b110x0x10x0x0x11: bits_out=15'b110101101010111;
        15'b10x10x10x0x0x11: bits_out=15'b101101101010111;
        15'b0x110x10x0x0x11: bits_out=15'b011101101010111;
        15'b11110x10x0x0x11: bits_out=15'b111101101010111;
        15'b10x0x110x0x0x11: bits_out=15'b101011101010111;
        15'b0x10x110x0x0x11: bits_out=15'b011011101010111;
        15'b1110x110x0x0x11: bits_out=15'b111011101010111;
        15'b0x0x1110x0x0x11: bits_out=15'b010111101010111;
        15'b110x1110x0x0x11: bits_out=15'b110111101010111;
        15'b10x11110x0x0x11: bits_out=15'b101111101010111;
        15'b0x111110x0x0x11: bits_out=15'b011111101010111;
        15'b11111110x0x0x11: bits_out=15'b111111101010111;
        15'b0x0x0x0x10x0x11: bits_out=15'b010101011010111;
        15'b110x0x0x10x0x11: bits_out=15'b110101011010111;
        15'b10x10x0x10x0x11: bits_out=15'b101101011010111;
        15'b0x110x0x10x0x11: bits_out=15'b011101011010111;
        15'b11110x0x10x0x11: bits_out=15'b111101011010111;
        15'b10x0x10x10x0x11: bits_out=15'b101011011010111;
        15'b0x10x10x10x0x11: bits_out=15'b011011011010111;
        15'b1110x10x10x0x11: bits_out=15'b111011011010111;
        15'b0x0x110x10x0x11: bits_out=15'b010111011010111;
        15'b110x110x10x0x11: bits_out=15'b110111011010111;
        15'b10x1110x10x0x11: bits_out=15'b101111011010111;
        15'b0x11110x10x0x11: bits_out=15'b011111011010111;
        15'b1111110x10x0x11: bits_out=15'b111111011010111;
        15'b10x0x0x110x0x11: bits_out=15'b101010111010111;
        15'b0x10x0x110x0x11: bits_out=15'b011010111010111;
        15'b1110x0x110x0x11: bits_out=15'b111010111010111;
        15'b0x0x10x110x0x11: bits_out=15'b010110111010111;
        15'b110x10x110x0x11: bits_out=15'b110110111010111;
        15'b10x110x110x0x11: bits_out=15'b101110111010111;
        15'b0x1110x110x0x11: bits_out=15'b011110111010111;
        15'b111110x110x0x11: bits_out=15'b111110111010111;
        15'b0x0x0x1110x0x11: bits_out=15'b010101111010111;
        15'b110x0x1110x0x11: bits_out=15'b110101111010111;
        15'b10x10x1110x0x11: bits_out=15'b101101111010111;
        15'b0x110x1110x0x11: bits_out=15'b011101111010111;
        15'b11110x1110x0x11: bits_out=15'b111101111010111;
        15'b10x0x11110x0x11: bits_out=15'b101011111010111;
        15'b0x10x11110x0x11: bits_out=15'b011011111010111;
        15'b1110x11110x0x11: bits_out=15'b111011111010111;
        15'b0x0x111110x0x11: bits_out=15'b010111111010111;
        15'b110x111110x0x11: bits_out=15'b110111111010111;
        15'b10x1111110x0x11: bits_out=15'b101111111010111;
        15'b0x11111110x0x11: bits_out=15'b011111111010111;
        15'b1111111110x0x11: bits_out=15'b111111111010111;
        15'b0x0x0x0x0x10x11: bits_out=15'b010101010110111;
        15'b110x0x0x0x10x11: bits_out=15'b110101010110111;
        15'b10x10x0x0x10x11: bits_out=15'b101101010110111;
        15'b0x110x0x0x10x11: bits_out=15'b011101010110111;
        15'b11110x0x0x10x11: bits_out=15'b111101010110111;
        15'b10x0x10x0x10x11: bits_out=15'b101011010110111;
        15'b0x10x10x0x10x11: bits_out=15'b011011010110111;
        15'b1110x10x0x10x11: bits_out=15'b111011010110111;
        15'b0x0x110x0x10x11: bits_out=15'b010111010110111;
        15'b110x110x0x10x11: bits_out=15'b110111010110111;
        15'b10x1110x0x10x11: bits_out=15'b101111010110111;
        15'b0x11110x0x10x11: bits_out=15'b011111010110111;
        15'b1111110x0x10x11: bits_out=15'b111111010110111;
        15'b10x0x0x10x10x11: bits_out=15'b101010110110111;
        15'b0x10x0x10x10x11: bits_out=15'b011010110110111;
        15'b1110x0x10x10x11: bits_out=15'b111010110110111;
        15'b0x0x10x10x10x11: bits_out=15'b010110110110111;
        15'b110x10x10x10x11: bits_out=15'b110110110110111;
        15'b10x110x10x10x11: bits_out=15'b101110110110111;
        15'b0x1110x10x10x11: bits_out=15'b011110110110111;
        15'b111110x10x10x11: bits_out=15'b111110110110111;
        15'b0x0x0x110x10x11: bits_out=15'b010101110110111;
        15'b110x0x110x10x11: bits_out=15'b110101110110111;
        15'b10x10x110x10x11: bits_out=15'b101101110110111;
        15'b0x110x110x10x11: bits_out=15'b011101110110111;
        15'b11110x110x10x11: bits_out=15'b111101110110111;
        15'b10x0x1110x10x11: bits_out=15'b101011110110111;
        15'b0x10x1110x10x11: bits_out=15'b011011110110111;
        15'b1110x1110x10x11: bits_out=15'b111011110110111;
        15'b0x0x11110x10x11: bits_out=15'b010111110110111;
        15'b110x11110x10x11: bits_out=15'b110111110110111;
        15'b10x111110x10x11: bits_out=15'b101111110110111;
        15'b0x1111110x10x11: bits_out=15'b011111110110111;
        15'b111111110x10x11: bits_out=15'b111111110110111;
        15'b10x0x0x0x110x11: bits_out=15'b101010101110111;
        15'b0x10x0x0x110x11: bits_out=15'b011010101110111;
        15'b1110x0x0x110x11: bits_out=15'b111010101110111;
        15'b0x0x10x0x110x11: bits_out=15'b010110101110111;
        15'b110x10x0x110x11: bits_out=15'b110110101110111;
        15'b10x110x0x110x11: bits_out=15'b101110101110111;
        15'b0x1110x0x110x11: bits_out=15'b011110101110111;
        15'b111110x0x110x11: bits_out=15'b111110101110111;
        15'b0x0x0x10x110x11: bits_out=15'b010101101110111;
        15'b110x0x10x110x11: bits_out=15'b110101101110111;
        15'b10x10x10x110x11: bits_out=15'b101101101110111;
        15'b0x110x10x110x11: bits_out=15'b011101101110111;
        15'b11110x10x110x11: bits_out=15'b111101101110111;
        15'b10x0x110x110x11: bits_out=15'b101011101110111;
        15'b0x10x110x110x11: bits_out=15'b011011101110111;
        15'b1110x110x110x11: bits_out=15'b111011101110111;
        15'b0x0x1110x110x11: bits_out=15'b010111101110111;
        15'b110x1110x110x11: bits_out=15'b110111101110111;
        15'b10x11110x110x11: bits_out=15'b101111101110111;
        15'b0x111110x110x11: bits_out=15'b011111101110111;
        15'b11111110x110x11: bits_out=15'b111111101110111;
        15'b0x0x0x0x1110x11: bits_out=15'b010101011110111;
        15'b110x0x0x1110x11: bits_out=15'b110101011110111;
        15'b10x10x0x1110x11: bits_out=15'b101101011110111;
        15'b0x110x0x1110x11: bits_out=15'b011101011110111;
        15'b11110x0x1110x11: bits_out=15'b111101011110111;
        15'b10x0x10x1110x11: bits_out=15'b101011011110111;
        15'b0x10x10x1110x11: bits_out=15'b011011011110111;
        15'b1110x10x1110x11: bits_out=15'b111011011110111;
        15'b0x0x110x1110x11: bits_out=15'b010111011110111;
        15'b110x110x1110x11: bits_out=15'b110111011110111;
        15'b10x1110x1110x11: bits_out=15'b101111011110111;
        15'b0x11110x1110x11: bits_out=15'b011111011110111;
        15'b1111110x1110x11: bits_out=15'b111111011110111;
        15'b10x0x0x11110x11: bits_out=15'b101010111110111;
        15'b0x10x0x11110x11: bits_out=15'b011010111110111;
        15'b1110x0x11110x11: bits_out=15'b111010111110111;
        15'b0x0x10x11110x11: bits_out=15'b010110111110111;
        15'b110x10x11110x11: bits_out=15'b110110111110111;
        15'b10x110x11110x11: bits_out=15'b101110111110111;
        15'b0x1110x11110x11: bits_out=15'b011110111110111;
        15'b111110x11110x11: bits_out=15'b111110111110111;
        15'b0x0x0x111110x11: bits_out=15'b010101111110111;
        15'b110x0x111110x11: bits_out=15'b110101111110111;
        15'b10x10x111110x11: bits_out=15'b101101111110111;
        15'b0x110x111110x11: bits_out=15'b011101111110111;
        15'b11110x111110x11: bits_out=15'b111101111110111;
        15'b10x0x1111110x11: bits_out=15'b101011111110111;
        15'b0x10x1111110x11: bits_out=15'b011011111110111;
        15'b1110x1111110x11: bits_out=15'b111011111110111;
        15'b0x0x11111110x11: bits_out=15'b010111111110111;
        15'b110x11111110x11: bits_out=15'b110111111110111;
        15'b10x111111110x11: bits_out=15'b101111111110111;
        15'b0x1111111110x11: bits_out=15'b011111111110111;
        15'b111111111110x11: bits_out=15'b111111111110111;
        15'b0x0x0x0x0x0x111: bits_out=15'b010101010101111;
        15'b110x0x0x0x0x111: bits_out=15'b110101010101111;
        15'b10x10x0x0x0x111: bits_out=15'b101101010101111;
        15'b0x110x0x0x0x111: bits_out=15'b011101010101111;
        15'b11110x0x0x0x111: bits_out=15'b111101010101111;
        15'b10x0x10x0x0x111: bits_out=15'b101011010101111;
        15'b0x10x10x0x0x111: bits_out=15'b011011010101111;
        15'b1110x10x0x0x111: bits_out=15'b111011010101111;
        15'b0x0x110x0x0x111: bits_out=15'b010111010101111;
        15'b110x110x0x0x111: bits_out=15'b110111010101111;
        15'b10x1110x0x0x111: bits_out=15'b101111010101111;
        15'b0x11110x0x0x111: bits_out=15'b011111010101111;
        15'b1111110x0x0x111: bits_out=15'b111111010101111;
        15'b10x0x0x10x0x111: bits_out=15'b101010110101111;
        15'b0x10x0x10x0x111: bits_out=15'b011010110101111;
        15'b1110x0x10x0x111: bits_out=15'b111010110101111;
        15'b0x0x10x10x0x111: bits_out=15'b010110110101111;
        15'b110x10x10x0x111: bits_out=15'b110110110101111;
        15'b10x110x10x0x111: bits_out=15'b101110110101111;
        15'b0x1110x10x0x111: bits_out=15'b011110110101111;
        15'b111110x10x0x111: bits_out=15'b111110110101111;
        15'b0x0x0x110x0x111: bits_out=15'b010101110101111;
        15'b110x0x110x0x111: bits_out=15'b110101110101111;
        15'b10x10x110x0x111: bits_out=15'b101101110101111;
        15'b0x110x110x0x111: bits_out=15'b011101110101111;
        15'b11110x110x0x111: bits_out=15'b111101110101111;
        15'b10x0x1110x0x111: bits_out=15'b101011110101111;
        15'b0x10x1110x0x111: bits_out=15'b011011110101111;
        15'b1110x1110x0x111: bits_out=15'b111011110101111;
        15'b0x0x11110x0x111: bits_out=15'b010111110101111;
        15'b110x11110x0x111: bits_out=15'b110111110101111;
        15'b10x111110x0x111: bits_out=15'b101111110101111;
        15'b0x1111110x0x111: bits_out=15'b011111110101111;
        15'b111111110x0x111: bits_out=15'b111111110101111;
        15'b10x0x0x0x10x111: bits_out=15'b101010101101111;
        15'b0x10x0x0x10x111: bits_out=15'b011010101101111;
        15'b1110x0x0x10x111: bits_out=15'b111010101101111;
        15'b0x0x10x0x10x111: bits_out=15'b010110101101111;
        15'b110x10x0x10x111: bits_out=15'b110110101101111;
        15'b10x110x0x10x111: bits_out=15'b101110101101111;
        15'b0x1110x0x10x111: bits_out=15'b011110101101111;
        15'b111110x0x10x111: bits_out=15'b111110101101111;
        15'b0x0x0x10x10x111: bits_out=15'b010101101101111;
        15'b110x0x10x10x111: bits_out=15'b110101101101111;
        15'b10x10x10x10x111: bits_out=15'b101101101101111;
        15'b0x110x10x10x111: bits_out=15'b011101101101111;
        15'b11110x10x10x111: bits_out=15'b111101101101111;
        15'b10x0x110x10x111: bits_out=15'b101011101101111;
        15'b0x10x110x10x111: bits_out=15'b011011101101111;
        15'b1110x110x10x111: bits_out=15'b111011101101111;
        15'b0x0x1110x10x111: bits_out=15'b010111101101111;
        15'b110x1110x10x111: bits_out=15'b110111101101111;
        15'b10x11110x10x111: bits_out=15'b101111101101111;
        15'b0x111110x10x111: bits_out=15'b011111101101111;
        15'b11111110x10x111: bits_out=15'b111111101101111;
        15'b0x0x0x0x110x111: bits_out=15'b010101011101111;
        15'b110x0x0x110x111: bits_out=15'b110101011101111;
        15'b10x10x0x110x111: bits_out=15'b101101011101111;
        15'b0x110x0x110x111: bits_out=15'b011101011101111;
        15'b11110x0x110x111: bits_out=15'b111101011101111;
        15'b10x0x10x110x111: bits_out=15'b101011011101111;
        15'b0x10x10x110x111: bits_out=15'b011011011101111;
        15'b1110x10x110x111: bits_out=15'b111011011101111;
        15'b0x0x110x110x111: bits_out=15'b010111011101111;
        15'b110x110x110x111: bits_out=15'b110111011101111;
        15'b10x1110x110x111: bits_out=15'b101111011101111;
        15'b0x11110x110x111: bits_out=15'b011111011101111;
        15'b1111110x110x111: bits_out=15'b111111011101111;
        15'b10x0x0x1110x111: bits_out=15'b101010111101111;
        15'b0x10x0x1110x111: bits_out=15'b011010111101111;
        15'b1110x0x1110x111: bits_out=15'b111010111101111;
        15'b0x0x10x1110x111: bits_out=15'b010110111101111;
        15'b110x10x1110x111: bits_out=15'b110110111101111;
        15'b10x110x1110x111: bits_out=15'b101110111101111;
        15'b0x1110x1110x111: bits_out=15'b011110111101111;
        15'b111110x1110x111: bits_out=15'b111110111101111;
        15'b0x0x0x11110x111: bits_out=15'b010101111101111;
        15'b110x0x11110x111: bits_out=15'b110101111101111;
        15'b10x10x11110x111: bits_out=15'b101101111101111;
        15'b0x110x11110x111: bits_out=15'b011101111101111;
        15'b11110x11110x111: bits_out=15'b111101111101111;
        15'b10x0x111110x111: bits_out=15'b101011111101111;
        15'b0x10x111110x111: bits_out=15'b011011111101111;
        15'b1110x111110x111: bits_out=15'b111011111101111;
        15'b0x0x1111110x111: bits_out=15'b010111111101111;
        15'b110x1111110x111: bits_out=15'b110111111101111;
        15'b10x11111110x111: bits_out=15'b101111111101111;
        15'b0x111111110x111: bits_out=15'b011111111101111;
        15'b11111111110x111: bits_out=15'b111111111101111;
        15'b10x0x0x0x0x1111: bits_out=15'b101010101011111;
        15'b0x10x0x0x0x1111: bits_out=15'b011010101011111;
        15'b1110x0x0x0x1111: bits_out=15'b111010101011111;
        15'b0x0x10x0x0x1111: bits_out=15'b010110101011111;
        15'b110x10x0x0x1111: bits_out=15'b110110101011111;
        15'b10x110x0x0x1111: bits_out=15'b101110101011111;
        15'b0x1110x0x0x1111: bits_out=15'b011110101011111;
        15'b111110x0x0x1111: bits_out=15'b111110101011111;
        15'b0x0x0x10x0x1111: bits_out=15'b010101101011111;
        15'b110x0x10x0x1111: bits_out=15'b110101101011111;
        15'b10x10x10x0x1111: bits_out=15'b101101101011111;
        15'b0x110x10x0x1111: bits_out=15'b011101101011111;
        15'b11110x10x0x1111: bits_out=15'b111101101011111;
        15'b10x0x110x0x1111: bits_out=15'b101011101011111;
        15'b0x10x110x0x1111: bits_out=15'b011011101011111;
        15'b1110x110x0x1111: bits_out=15'b111011101011111;
        15'b0x0x1110x0x1111: bits_out=15'b010111101011111;
        15'b110x1110x0x1111: bits_out=15'b110111101011111;
        15'b10x11110x0x1111: bits_out=15'b101111101011111;
        15'b0x111110x0x1111: bits_out=15'b011111101011111;
        15'b11111110x0x1111: bits_out=15'b111111101011111;
        15'b0x0x0x0x10x1111: bits_out=15'b010101011011111;
        15'b110x0x0x10x1111: bits_out=15'b110101011011111;
        15'b10x10x0x10x1111: bits_out=15'b101101011011111;
        15'b0x110x0x10x1111: bits_out=15'b011101011011111;
        15'b11110x0x10x1111: bits_out=15'b111101011011111;
        15'b10x0x10x10x1111: bits_out=15'b101011011011111;
        15'b0x10x10x10x1111: bits_out=15'b011011011011111;
        15'b1110x10x10x1111: bits_out=15'b111011011011111;
        15'b0x0x110x10x1111: bits_out=15'b010111011011111;
        15'b110x110x10x1111: bits_out=15'b110111011011111;
        15'b10x1110x10x1111: bits_out=15'b101111011011111;
        15'b0x11110x10x1111: bits_out=15'b011111011011111;
        15'b1111110x10x1111: bits_out=15'b111111011011111;
        15'b10x0x0x110x1111: bits_out=15'b101010111011111;
        15'b0x10x0x110x1111: bits_out=15'b011010111011111;
        15'b1110x0x110x1111: bits_out=15'b111010111011111;
        15'b0x0x10x110x1111: bits_out=15'b010110111011111;
        15'b110x10x110x1111: bits_out=15'b110110111011111;
        15'b10x110x110x1111: bits_out=15'b101110111011111;
        15'b0x1110x110x1111: bits_out=15'b011110111011111;
        15'b111110x110x1111: bits_out=15'b111110111011111;
        15'b0x0x0x1110x1111: bits_out=15'b010101111011111;
        15'b110x0x1110x1111: bits_out=15'b110101111011111;
        15'b10x10x1110x1111: bits_out=15'b101101111011111;
        15'b0x110x1110x1111: bits_out=15'b011101111011111;
        15'b11110x1110x1111: bits_out=15'b111101111011111;
        15'b10x0x11110x1111: bits_out=15'b101011111011111;
        15'b0x10x11110x1111: bits_out=15'b011011111011111;
        15'b1110x11110x1111: bits_out=15'b111011111011111;
        15'b0x0x111110x1111: bits_out=15'b010111111011111;
        15'b110x111110x1111: bits_out=15'b110111111011111;
        15'b10x1111110x1111: bits_out=15'b101111111011111;
        15'b0x11111110x1111: bits_out=15'b011111111011111;
        15'b1111111110x1111: bits_out=15'b111111111011111;
        15'b0x0x0x0x0x11111: bits_out=15'b010101010111111;
        15'b110x0x0x0x11111: bits_out=15'b110101010111111;
        15'b10x10x0x0x11111: bits_out=15'b101101010111111;
        15'b0x110x0x0x11111: bits_out=15'b011101010111111;
        15'b11110x0x0x11111: bits_out=15'b111101010111111;
        15'b10x0x10x0x11111: bits_out=15'b101011010111111;
        15'b0x10x10x0x11111: bits_out=15'b011011010111111;
        15'b1110x10x0x11111: bits_out=15'b111011010111111;
        15'b0x0x110x0x11111: bits_out=15'b010111010111111;
        15'b110x110x0x11111: bits_out=15'b110111010111111;
        15'b10x1110x0x11111: bits_out=15'b101111010111111;
        15'b0x11110x0x11111: bits_out=15'b011111010111111;
        15'b1111110x0x11111: bits_out=15'b111111010111111;
        15'b10x0x0x10x11111: bits_out=15'b101010110111111;
        15'b0x10x0x10x11111: bits_out=15'b011010110111111;
        15'b1110x0x10x11111: bits_out=15'b111010110111111;
        15'b0x0x10x10x11111: bits_out=15'b010110110111111;
        15'b110x10x10x11111: bits_out=15'b110110110111111;
        15'b10x110x10x11111: bits_out=15'b101110110111111;
        15'b0x1110x10x11111: bits_out=15'b011110110111111;
        15'b111110x10x11111: bits_out=15'b111110110111111;
        15'b0x0x0x110x11111: bits_out=15'b010101110111111;
        15'b110x0x110x11111: bits_out=15'b110101110111111;
        15'b10x10x110x11111: bits_out=15'b101101110111111;
        15'b0x110x110x11111: bits_out=15'b011101110111111;
        15'b11110x110x11111: bits_out=15'b111101110111111;
        15'b10x0x1110x11111: bits_out=15'b101011110111111;
        15'b0x10x1110x11111: bits_out=15'b011011110111111;
        15'b1110x1110x11111: bits_out=15'b111011110111111;
        15'b0x0x11110x11111: bits_out=15'b010111110111111;
        15'b110x11110x11111: bits_out=15'b110111110111111;
        15'b10x111110x11111: bits_out=15'b101111110111111;
        15'b0x1111110x11111: bits_out=15'b011111110111111;
        15'b111111110x11111: bits_out=15'b111111110111111;
        15'b10x0x0x0x111111: bits_out=15'b101010101111111;
        15'b0x10x0x0x111111: bits_out=15'b011010101111111;
        15'b1110x0x0x111111: bits_out=15'b111010101111111;
        15'b0x0x10x0x111111: bits_out=15'b010110101111111;
        15'b110x10x0x111111: bits_out=15'b110110101111111;
        15'b10x110x0x111111: bits_out=15'b101110101111111;
        15'b0x1110x0x111111: bits_out=15'b011110101111111;
        15'b111110x0x111111: bits_out=15'b111110101111111;
        15'b0x0x0x10x111111: bits_out=15'b010101101111111;
        15'b110x0x10x111111: bits_out=15'b110101101111111;
        15'b10x10x10x111111: bits_out=15'b101101101111111;
        15'b0x110x10x111111: bits_out=15'b011101101111111;
        15'b11110x10x111111: bits_out=15'b111101101111111;
        15'b10x0x110x111111: bits_out=15'b101011101111111;
        15'b0x10x110x111111: bits_out=15'b011011101111111;
        15'b1110x110x111111: bits_out=15'b111011101111111;
        15'b0x0x1110x111111: bits_out=15'b010111101111111;
        15'b110x1110x111111: bits_out=15'b110111101111111;
        15'b10x11110x111111: bits_out=15'b101111101111111;
        15'b0x111110x111111: bits_out=15'b011111101111111;
        15'b11111110x111111: bits_out=15'b111111101111111;
        15'b0x0x0x0x1111111: bits_out=15'b010101011111111;
        15'b110x0x0x1111111: bits_out=15'b110101011111111;
        15'b10x10x0x1111111: bits_out=15'b101101011111111;
        15'b0x110x0x1111111: bits_out=15'b011101011111111;
        15'b11110x0x1111111: bits_out=15'b111101011111111;
        15'b10x0x10x1111111: bits_out=15'b101011011111111;
        15'b0x10x10x1111111: bits_out=15'b011011011111111;
        15'b1110x10x1111111: bits_out=15'b111011011111111;
        15'b0x0x110x1111111: bits_out=15'b010111011111111;
        15'b110x110x1111111: bits_out=15'b110111011111111;
        15'b10x1110x1111111: bits_out=15'b101111011111111;
        15'b0x11110x1111111: bits_out=15'b011111011111111;
        15'b1111110x1111111: bits_out=15'b111111011111111;
        15'b10x0x0x11111111: bits_out=15'b101010111111111;
        15'b0x10x0x11111111: bits_out=15'b011010111111111;
        15'b1110x0x11111111: bits_out=15'b111010111111111;
        15'b0x0x10x11111111: bits_out=15'b010110111111111;
        15'b110x10x11111111: bits_out=15'b110110111111111;
        15'b10x110x11111111: bits_out=15'b101110111111111;
        15'b0x1110x11111111: bits_out=15'b011110111111111;
        15'b111110x11111111: bits_out=15'b111110111111111;
        15'b0x0x0x111111111: bits_out=15'b010101111111111;
        15'b110x0x111111111: bits_out=15'b110101111111111;
        15'b10x10x111111111: bits_out=15'b101101111111111;
        15'b0x110x111111111: bits_out=15'b011101111111111;
        15'b11110x111111111: bits_out=15'b111101111111111;
        15'b10x0x1111111111: bits_out=15'b101011111111111;
        15'b0x10x1111111111: bits_out=15'b011011111111111;
        15'b1110x1111111111: bits_out=15'b111011111111111;
        15'b0x0x11111111111: bits_out=15'b010111111111111;
        15'b110x11111111111: bits_out=15'b110111111111111;
        15'b10x111111111111: bits_out=15'b101111111111111;
        15'b0x1111111111111: bits_out=15'b011111111111111;
        15'b111111111111111: bits_out=15'b111111111111111;
    endcase
  end
endmodule
