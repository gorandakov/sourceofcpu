/*
Copyright 2022 Goran Dakov

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

module fpucadd_compress(clk,R,C,A_out,B_out,or1,and1);
  input clk;
  input [64:0] R;
  input [64:0] C;
  output [127:0] A_out;
  output [127:0] B_out;
  input or1;
  input and1;//and1 inverse of or1
  reg REGS_0;
  reg REGS_1;
  reg REGS_2;
  reg REGS_3;
  reg REGS_4;
  reg REGS_5;
  reg REGS_6;
  reg REGS_7;
  reg REGS_8;
  reg REGS_9;
  reg REGS_10;
  reg REGS_11;
  reg REGS_12;
  reg REGS_13;
  reg REGS_14;
  reg REGS_15;
  reg REGS_16;
  reg REGS_17;
  reg REGS_18;
  reg REGS_19;
  reg REGS_20;
  reg REGS_21;
  reg REGS_22;
  reg REGS_23;
  reg REGS_24;
  reg REGS_25;
  reg REGS_26;
  reg REGS_27;
  reg REGS_28;
  reg REGS_29;
  reg REGS_30;
  reg REGS_31;
  reg REGS_32;
  reg REGS_33;
  reg REGS_34;
  reg REGS_35;
  reg REGS_36;
  reg REGS_37;
  reg REGS_38;
  reg REGS_39;
  reg REGS_40;
  reg REGS_41;
  reg REGS_42;
  reg REGS_43;
  reg REGS_44;
  reg REGS_45;
  reg REGS_46;
  reg REGS_47;
  reg REGS_48;
  reg REGS_49;
  reg REGS_50;
  reg REGS_51;
  reg REGS_52;
  reg REGS_53;
  reg REGS_54;
  reg REGS_55;
  reg REGS_56;
  reg REGS_57;
  reg REGS_58;
  reg REGS_59;
  reg REGS_60;
  reg REGS_61;
  reg REGS_62;
  reg REGS_63;
  reg REGS_64;
  reg REGS_65;
  reg REGS_66;
  reg REGS_67;
  reg REGS_68;
  reg REGS_69;
  reg REGS_70;
  reg REGS_71;
  reg REGS_72;
  reg REGS_73;
  reg REGS_74;
  reg REGS_75;
  reg REGS_76;
  reg REGS_77;
  reg REGS_78;
  reg REGS_79;
  reg REGS_80;
  reg REGS_81;
  reg REGS_82;
  reg REGS_83;
  reg REGS_84;
  reg REGS_85;
  reg REGS_86;
  reg REGS_87;
  reg REGS_88;
  reg REGS_89;
  reg REGS_90;
  reg REGS_91;
  reg REGS_92;
  reg REGS_93;
  reg REGS_94;
  reg REGS_95;
  reg REGS_96;
  reg REGS_97;
  reg REGS_98;
  reg REGS_99;
  reg REGS_100;
  reg REGS_101;
  reg REGS_102;
  reg REGS_103;
  reg REGS_104;
  reg REGS_105;
  reg REGS_106;
  reg REGS_107;
  reg REGS_108;
  reg REGS_109;
  reg REGS_110;
  reg REGS_111;
  reg REGS_112;
  reg REGS_113;
  reg REGS_114;
  reg REGS_115;
  reg REGS_116;
  reg REGS_117;
  reg REGS_118;
  reg REGS_119;
  reg REGS_120;
  reg REGS_121;
  reg REGS_122;
  reg REGS_123;
  reg REGS_124;
  reg REGS_125;
  reg REGS_126;
  reg REGS_127;
  reg REGS_128;
  reg REGS_129;
  reg REGS_130;
  reg REGS_131;
  reg REGS_132;
  reg REGS_133;
  reg REGS_134;
  reg REGS_135;
  reg REGS_136;
  reg REGS_137;
  reg REGS_138;
  reg REGS_139;
  reg REGS_140;
  reg REGS_141;
  reg REGS_142;
  reg REGS_143;
  reg REGS_144;
  reg REGS_145;
  reg REGS_146;
  reg REGS_147;
  reg REGS_148;
  reg REGS_149;
  reg REGS_150;
  reg REGS_151;
  reg REGS_152;
  reg REGS_153;
  reg REGS_154;
  reg REGS_155;
  reg REGS_156;
  reg REGS_157;
  reg REGS_158;
  reg REGS_159;
  reg REGS_160;
  reg REGS_161;
  reg REGS_162;
  reg REGS_163;
  reg REGS_164;
  reg REGS_165;
  reg REGS_166;
  reg REGS_167;
  reg REGS_168;
  reg REGS_169;
  reg REGS_170;
  reg REGS_171;
  reg REGS_172;
  reg REGS_173;
  reg REGS_174;
  reg REGS_175;
  reg REGS_176;
  reg REGS_177;
  reg REGS_178;
  reg REGS_179;
  reg REGS_180;
  reg REGS_181;
  reg REGS_182;
  reg REGS_183;
  reg REGS_184;
  reg REGS_185;
  reg REGS_186;
  reg REGS_187;
  reg REGS_188;
  reg REGS_189;
  reg REGS_190;
  reg REGS_191;
  reg REGS_192;
  reg REGS_193;
  reg REGS_194;
  reg REGS_195;
  reg REGS_196;
  reg REGS_197;
  reg REGS_198;
  reg REGS_199;
  reg REGS_200;
  reg REGS_201;
  reg REGS_202;
  reg REGS_203;
  reg REGS_204;
  reg REGS_205;
  reg REGS_206;
  reg REGS_207;
  reg REGS_208;
  reg REGS_209;
  reg REGS_210;
  reg REGS_211;
  reg REGS_212;
  reg REGS_213;
  reg REGS_214;
  reg REGS_215;
  reg REGS_216;
  reg REGS_217;
  reg REGS_218;
  reg REGS_219;
  reg REGS_220;
  reg REGS_221;
  reg REGS_222;
  reg REGS_223;
  reg REGS_224;
  reg REGS_225;
  reg REGS_226;
  reg REGS_227;
  reg REGS_228;
  reg REGS_229;
  reg REGS_230;
  reg REGS_231;
  reg REGS_232;
  reg REGS_233;
  reg REGS_234;
  reg REGS_235;
  reg REGS_236;
  reg REGS_237;
  reg REGS_238;
  reg REGS_239;
  reg REGS_240;
  reg REGS_241;
  reg REGS_242;
  reg REGS_243;
  reg REGS_244;
  reg REGS_245;
  reg REGS_246;
  reg REGS_247;
  reg REGS_248;
  reg REGS_249;
  reg REGS_250;
  reg REGS_251;
  reg REGS_252;
  reg REGS_253;
  reg REGS_254;
  reg REGS_255;
  reg REGS_256;
  reg REGS_257;
  reg REGS_258;
  reg REGS_259;
  reg REGS_260;
  reg REGS_261;
  reg REGS_262;
  reg REGS_263;
  reg REGS_264;
  reg REGS_265;
  reg REGS_266;
  reg REGS_267;
  reg REGS_268;
  reg REGS_269;
  reg REGS_270;
  reg REGS_271;
  reg REGS_272;
  reg REGS_273;
  reg REGS_274;
  reg REGS_275;
  reg REGS_276;
  reg REGS_277;
  reg REGS_278;
  reg REGS_279;
  reg REGS_280;
  reg REGS_281;
  reg REGS_282;
  reg REGS_283;
  reg REGS_284;
  reg REGS_285;
  reg REGS_286;
  reg REGS_287;
  reg REGS_288;
  reg REGS_289;
  reg REGS_290;
  reg REGS_291;
  reg REGS_292;
  reg REGS_293;
  reg REGS_294;
  reg REGS_295;
  reg REGS_296;
  reg REGS_297;
  reg REGS_298;
  reg REGS_299;
  reg REGS_300;
  reg REGS_301;
  reg REGS_302;
  reg REGS_303;
  reg REGS_304;
  reg REGS_305;
  reg REGS_306;
  reg REGS_307;
  reg REGS_308;
  reg REGS_309;
  reg REGS_310;
  reg REGS_311;
  reg REGS_312;
  reg REGS_313;
  reg REGS_314;
  reg REGS_315;
  reg REGS_316;
  reg REGS_317;
  reg REGS_318;
  reg REGS_319;
  reg REGS_320;
  reg REGS_321;
  reg REGS_322;
  reg REGS_323;
  reg REGS_324;
  reg REGS_325;
  reg REGS_326;
  reg REGS_327;
  reg REGS_328;
  reg REGS_329;
  reg REGS_330;
  reg REGS_331;
  reg REGS_332;
  reg REGS_333;
  reg REGS_334;
  reg REGS_335;
  reg REGS_336;
  reg REGS_337;
  reg REGS_338;
  reg REGS_339;
  reg REGS_340;
  reg REGS_341;
  reg REGS_342;
  reg REGS_343;
  reg REGS_344;
  reg REGS_345;
  reg REGS_346;
  reg REGS_347;
  reg REGS_348;
  reg REGS_349;
  reg REGS_350;
  reg REGS_351;
  reg REGS_352;
  reg REGS_353;
  reg REGS_354;
  reg REGS_355;
  reg REGS_356;
  reg REGS_357;
  reg REGS_358;
  reg REGS_359;
  reg REGS_360;
  reg REGS_361;
  reg REGS_362;
  reg REGS_363;
  reg REGS_364;
  reg REGS_365;
  reg REGS_366;
  reg REGS_367;
  reg REGS_368;
  reg REGS_369;
  reg REGS_370;
  reg REGS_371;
  reg REGS_372;
  reg REGS_373;
  reg REGS_374;
  reg REGS_375;
  reg REGS_376;
  reg REGS_377;
  reg REGS_378;
  reg REGS_379;
  reg REGS_380;
  reg REGS_381;
  reg REGS_382;
  reg REGS_383;
  reg REGS_384;
  reg REGS_385;
  reg REGS_386;
  reg REGS_387;
  reg REGS_388;
  reg REGS_389;
  reg REGS_390;
  reg REGS_391;
  reg REGS_392;
  reg REGS_393;
  reg REGS_394;
  reg REGS_395;
  reg REGS_396;
  reg REGS_397;
  reg REGS_398;
  reg REGS_399;
  reg REGS_400;
  reg REGS_401;
  reg REGS_402;
  reg REGS_403;
  reg REGS_404;
  reg REGS_405;
  reg REGS_406;
  reg REGS_407;
  reg REGS_408;
  reg REGS_409;
  reg REGS_410;
  reg REGS_411;
  reg REGS_412;
  reg REGS_413;
  reg REGS_414;
  reg REGS_415;
  reg REGS_416;
  reg REGS_417;
  reg REGS_418;
  reg REGS_419;
  reg REGS_420;
  reg REGS_421;
  reg REGS_422;
  reg REGS_423;
  reg REGS_424;
  reg REGS_425;
  reg REGS_426;
  reg REGS_427;
  reg REGS_428;
  reg REGS_429;
  reg REGS_430;
  reg REGS_431;
  reg REGS_432;
  reg REGS_433;
  reg REGS_434;
  reg REGS_435;
  reg REGS_436;
  reg REGS_437;
  reg REGS_438;
  reg REGS_439;
  reg REGS_440;
  reg REGS_441;
  reg REGS_442;
  reg REGS_443;
  reg REGS_444;
  reg REGS_445;
  reg REGS_446;
  reg REGS_447;
  reg REGS_448;
  reg REGS_449;
  reg REGS_450;
  reg REGS_451;
  reg REGS_452;
  reg REGS_453;
  reg REGS_454;
  reg REGS_455;
  reg REGS_456;
  reg REGS_457;
  reg REGS_458;
  reg REGS_459;
  reg REGS_460;
  reg REGS_461;
  reg REGS_462;
  reg REGS_463;
  reg REGS_464;
  reg REGS_465;
  reg REGS_466;
  reg REGS_467;
  reg REGS_468;
  reg REGS_469;
  reg REGS_470;
  reg REGS_471;
  reg REGS_472;
  reg REGS_473;
  reg REGS_474;
  reg REGS_475;
  reg REGS_476;
  reg REGS_477;
  reg REGS_478;
  reg REGS_479;
  reg REGS_480;
  reg REGS_481;
  reg REGS_482;
  reg REGS_483;
  reg REGS_484;
  reg REGS_485;
  reg REGS_486;
  reg REGS_487;
  reg REGS_488;
  reg REGS_489;
  reg REGS_490;
  reg REGS_491;
  reg REGS_492;
  reg REGS_493;
  reg REGS_494;
  reg REGS_495;
  reg REGS_496;
  reg REGS_497;
  reg REGS_498;
  reg REGS_499;
  reg REGS_500;
  reg REGS_501;
  reg REGS_502;
  reg REGS_503;
  reg REGS_504;
  reg REGS_505;
  reg REGS_506;
  reg REGS_507;
  reg REGS_508;
  reg REGS_509;
  reg REGS_510;
  reg REGS_511;
  reg REGS_512;
  reg REGS_513;
  reg REGS_514;
  reg REGS_515;
  reg REGS_516;
  reg REGS_517;
  reg REGS_518;
  reg REGS_519;
  reg REGS_520;
  reg REGS_521;
  reg REGS_522;
  reg REGS_523;
  reg REGS_524;
  reg REGS_525;
  reg REGS_526;
  reg REGS_527;
  reg REGS_528;
  reg REGS_529;
  reg REGS_530;
  reg REGS_531;
  reg REGS_532;
  reg REGS_533;
  reg REGS_534;
  reg REGS_535;
  reg REGS_536;
  reg REGS_537;
  reg REGS_538;
  reg REGS_539;
  reg REGS_540;
  reg REGS_541;
  reg REGS_542;
  reg REGS_543;
  reg REGS_544;
  reg REGS_545;
  reg REGS_546;
  reg REGS_547;
  reg REGS_548;
  reg REGS_549;
  reg REGS_550;
  reg REGS_551;
  reg REGS_552;
  reg REGS_553;
  reg REGS_554;
  reg REGS_555;
  reg REGS_556;
  reg REGS_557;
  reg REGS_558;
  reg REGS_559;
  reg REGS_560;
  reg REGS_561;
  reg REGS_562;
  reg REGS_563;
  reg REGS_564;
  reg REGS_565;
  reg REGS_566;
  reg REGS_567;
  reg REGS_568;
  reg REGS_569;
  reg REGS_570;
  reg REGS_571;
  reg REGS_572;
  reg REGS_573;
  reg REGS_574;
  reg REGS_575;
  reg REGS_576;
  reg REGS_577;
  reg REGS_578;
  reg REGS_579;
  reg REGS_580;
  reg REGS_581;
  reg REGS_582;
  reg REGS_583;
  reg REGS_584;
  reg REGS_585;
  reg REGS_586;
  reg REGS_587;
  reg REGS_588;
  reg REGS_589;
  reg REGS_590;
  reg REGS_591;
  reg REGS_592;
  reg REGS_593;
  reg REGS_594;
  reg REGS_595;
  reg REGS_596;
  reg REGS_597;
  reg REGS_598;
  reg REGS_599;
  reg REGS_600;
  reg REGS_601;
  reg REGS_602;
  reg REGS_603;
  reg REGS_604;
  reg REGS_605;
  reg REGS_606;
  reg REGS_607;
  reg REGS_608;
  reg REGS_609;
  reg REGS_610;
  reg REGS_611;
  reg REGS_612;
  reg REGS_613;
  reg REGS_614;
  reg REGS_615;
  reg REGS_616;
  reg REGS_617;
  reg REGS_618;
  reg REGS_619;
  reg REGS_620;
  reg REGS_621;
  reg REGS_622;
  reg REGS_623;
  reg REGS_624;
  reg REGS_625;
  reg REGS_626;
  reg REGS_627;
  reg REGS_628;
  reg REGS_629;
  reg REGS_630;
  reg REGS_631;
  reg REGS_632;
  reg REGS_633;
  reg REGS_634;
  reg REGS_635;
  reg REGS_636;
  reg REGS_637;
  reg REGS_638;
  reg REGS_639;
  reg REGS_640;
  reg REGS_641;
  reg REGS_642;
  reg REGS_643;
  reg REGS_644;
  reg REGS_645;
  reg REGS_646;
  reg REGS_647;
  reg REGS_648;
  reg REGS_649;
  reg REGS_650;
  reg REGS_651;
  reg REGS_652;
  reg REGS_653;
  reg REGS_654;
  reg REGS_655;
  reg REGS_656;
  reg REGS_657;
  reg REGS_658;
  reg REGS_659;
  reg REGS_660;
  reg REGS_661;
  reg REGS_662;
  reg REGS_663;
  reg REGS_664;
  reg REGS_665;
  reg REGS_666;
  reg REGS_667;
  reg REGS_668;
  reg REGS_669;
  reg REGS_670;
  reg REGS_671;
  reg REGS_672;
  reg REGS_673;
  reg REGS_674;
  reg REGS_675;
  reg REGS_676;
  reg REGS_677;
  reg REGS_678;
  reg REGS_679;
  reg REGS_680;
  reg REGS_681;
  reg REGS_682;
  reg REGS_683;
  reg REGS_684;
  reg REGS_685;
  reg REGS_686;
  reg REGS_687;
  reg REGS_688;
  reg REGS_689;
  reg REGS_690;
  reg REGS_691;
  reg REGS_692;
  reg REGS_693;
  reg REGS_694;
  reg REGS_695;
  reg REGS_696;
  reg REGS_697;
  reg REGS_698;
  reg REGS_699;
  reg REGS_700;
  reg REGS_701;
  reg REGS_702;
  reg REGS_703;
  reg REGS_704;
  reg REGS_705;
  reg REGS_706;
  reg REGS_707;
  reg REGS_708;
  reg REGS_709;
  reg REGS_710;
  reg REGS_711;
  reg REGS_712;
  reg REGS_713;
  reg REGS_714;
  reg REGS_715;
  reg REGS_716;
  reg REGS_717;
  reg REGS_718;
  reg REGS_719;
  reg REGS_720;
  reg REGS_721;
  reg REGS_722;
  reg REGS_723;
  reg REGS_724;
  reg REGS_725;
  reg REGS_726;
  reg REGS_727;
  reg REGS_728;
  reg REGS_729;
  reg REGS_730;
  reg REGS_731;
  reg REGS_732;
  reg REGS_733;
  reg REGS_734;
  reg REGS_735;
  reg REGS_736;
  reg REGS_737;
  reg REGS_738;
  reg REGS_739;
  reg REGS_740;
  reg REGS_741;
  reg REGS_742;
  reg REGS_743;
  reg REGS_744;
  reg REGS_745;
  reg REGS_746;
  reg REGS_747;
  reg REGS_748;
  reg REGS_749;
  reg REGS_750;
  reg REGS_751;
  reg REGS_752;
  reg REGS_753;
  reg REGS_754;
  reg REGS_755;
  reg REGS_756;
  reg REGS_757;
  reg REGS_758;
  reg REGS_759;
  reg REGS_760;
  reg REGS_761;
  reg REGS_762;
  reg REGS_763;
  reg REGS_764;
  reg REGS_765;
  reg REGS_766;
  reg REGS_767;
  reg REGS_768;
  reg REGS_769;
  reg REGS_770;
  reg REGS_771;
  reg REGS_772;
  reg REGS_773;
  reg REGS_774;
  reg REGS_775;
  reg REGS_776;
  reg REGS_777;
  reg REGS_778;
  reg REGS_779;
  reg REGS_780;
  reg REGS_781;
  reg REGS_782;
  reg REGS_783;
  reg REGS_784;
  reg REGS_785;
  reg REGS_786;
  reg REGS_787;
  reg REGS_788;
  reg REGS_789;
  reg REGS_790;
  reg REGS_791;
  reg REGS_792;
  reg REGS_793;
  reg REGS_794;
  reg REGS_795;
  reg REGS_796;
  reg REGS_797;
  reg REGS_798;
  reg REGS_799;
  reg REGS_800;
  reg REGS_801;
  reg REGS_802;
  reg REGS_803;
  reg REGS_804;
  reg REGS_805;
  reg REGS_806;
  reg REGS_807;
  reg REGS_808;
  reg REGS_809;
  reg REGS_810;
  reg REGS_811;
  reg REGS_812;
  reg REGS_813;
  reg REGS_814;
  reg REGS_815;
  reg REGS_816;
  reg REGS_817;
  reg REGS_818;
  reg REGS_819;
  reg REGS_820;
  reg REGS_821;
  reg REGS_822;
  reg REGS_823;
  reg REGS_824;
  reg REGS_825;
  reg REGS_826;
  reg REGS_827;
  reg REGS_828;
  reg REGS_829;
  reg REGS_830;
  reg REGS_831;
  reg REGS_832;
  reg REGS_833;
  reg REGS_834;
  reg REGS_835;
  reg REGS_836;
  reg REGS_837;
  reg REGS_838;
  reg REGS_839;
  reg REGS_840;
  reg REGS_841;
  reg REGS_842;
  reg REGS_843;
  reg REGS_844;
  reg REGS_845;
  reg REGS_846;
  reg REGS_847;
  reg REGS_848;
  reg REGS_849;
  reg REGS_850;
  reg REGS_851;
  reg REGS_852;
  reg REGS_853;
  reg REGS_854;
  reg REGS_855;
  reg REGS_856;
  reg REGS_857;
  reg REGS_858;
  reg REGS_859;
  reg REGS_860;
  reg REGS_861;
  reg REGS_862;
  reg REGS_863;
  reg REGS_864;
  reg REGS_865;
  reg REGS_866;
  reg REGS_867;
  reg REGS_868;
  reg REGS_869;
  reg REGS_870;
  reg REGS_871;
  reg REGS_872;
  reg REGS_873;
  reg REGS_874;
  reg REGS_875;
  reg REGS_876;
  reg REGS_877;
  reg REGS_878;
  reg REGS_879;
  reg REGS_880;
  reg REGS_881;
  reg REGS_882;
  reg REGS_883;
  reg REGS_884;
  reg REGS_885;
  reg REGS_886;
  reg REGS_887;
  reg REGS_888;
  reg REGS_889;
  reg REGS_890;
  reg REGS_891;
  reg REGS_892;
  reg REGS_893;
  reg REGS_894;
  reg REGS_895;
  reg REGS_896;
  reg REGS_897;
  reg REGS_898;
  reg REGS_899;
  reg REGS_900;
  reg REGS_901;
  reg REGS_902;
  reg REGS_903;
  reg REGS_904;
  reg REGS_905;
  reg REGS_906;
  reg REGS_907;
  reg REGS_908;
  reg REGS_909;
  reg REGS_910;
  reg REGS_911;
  reg REGS_912;
  reg REGS_913;
  reg REGS_914;
  reg REGS_915;
  reg REGS_916;
  reg REGS_917;
  reg REGS_918;
  reg REGS_919;
  reg REGS_920;
  reg REGS_921;
  reg REGS_922;
  reg REGS_923;
  reg REGS_924;
  reg REGS_925;
  reg REGS_926;
  reg REGS_927;
  reg REGS_928;
  reg REGS_929;
  reg REGS_930;
  reg REGS_931;
  reg REGS_932;
  reg REGS_933;
  reg REGS_934;
  reg REGS_935;
  reg REGS_936;
  reg REGS_937;
  reg REGS_938;
  reg REGS_939;
  reg REGS_940;
  reg REGS_941;
  reg REGS_942;
  reg REGS_943;
  reg REGS_944;
  reg REGS_945;
  reg REGS_946;
  reg REGS_947;
  reg REGS_948;
  reg REGS_949;
  reg REGS_950;
  reg REGS_951;
  reg REGS_952;
  reg REGS_953;
  reg REGS_954;
  reg REGS_955;
  reg REGS_956;
  reg REGS_957;
  reg REGS_958;
  reg REGS_959;
  reg REGS_960;
  reg REGS_961;
  reg REGS_962;
  reg REGS_963;
  reg REGS_964;
  reg REGS_965;
  reg REGS_966;
  reg REGS_967;
  reg REGS_968;
  reg REGS_969;
  reg REGS_970;
  reg REGS_971;
  reg REGS_972;
  reg REGS_973;
  reg REGS_974;
  reg REGS_975;
  reg REGS_976;
  reg REGS_977;
  reg REGS_978;
  reg REGS_979;
  reg REGS_980;
  reg REGS_981;
  reg REGS_982;
  reg REGS_983;
  reg REGS_984;
  reg REGS_985;
  reg REGS_986;
  reg REGS_987;
  reg REGS_988;
  reg REGS_989;
  reg REGS_990;
  reg REGS_991;
  reg REGS_992;
  reg REGS_993;
  reg REGS_994;
  reg REGS_995;
  reg REGS_996;
  reg REGS_997;
  reg REGS_998;
  reg REGS_999;
  reg REGS_1000;
  reg REGS_1001;
  reg REGS_1002;
  reg REGS_1003;
  reg REGS_1004;
  reg REGS_1005;
  reg REGS_1006;
  reg REGS_1007;
  reg REGS_1008;
  reg REGS_1009;
  reg REGS_1010;
  reg REGS_1011;
  reg REGS_1012;
  reg REGS_1013;
  reg REGS_1014;
  reg REGS_1015;
  reg REGS_1016;
  reg REGS_1017;
  reg REGS_1018;
  reg REGS_1019;
  reg REGS_1020;
  reg REGS_1021;
  reg REGS_1022;
  reg REGS_1023;
  reg REGS_1024;
  reg REGS_1025;
  reg REGS_1026;
  reg REGS_1027;
  reg REGS_1028;
  reg REGS_1029;
  reg REGS_1030;
  reg REGS_1031;
  reg REGS_1032;
  reg REGS_1033;
  reg REGS_1034;
  reg REGS_1035;
  reg REGS_1036;
  reg REGS_1037;
  reg REGS_1038;
  reg REGS_1039;
  reg REGS_1040;
  reg REGS_1041;
  reg REGS_1042;
  reg REGS_1043;
  reg REGS_1044;
  reg REGS_1045;
  reg REGS_1046;
  reg REGS_1047;
  reg REGS_1048;
  reg REGS_1049;
  reg REGS_1050;
  reg REGS_1051;
  reg REGS_1052;
  reg REGS_1053;
  reg REGS_1054;
  reg REGS_1055;
  reg REGS_1056;
  reg REGS_1057;
  reg REGS_1058;
  reg REGS_1059;
  reg REGS_1060;
  reg REGS_1061;
  reg REGS_1062;
  reg REGS_1063;
  reg REGS_1064;
  reg REGS_1065;
  reg REGS_1066;
  reg REGS_1067;
  reg REGS_1068;
  reg REGS_1069;
  reg REGS_1070;
  reg REGS_1071;
  reg REGS_1072;
  reg REGS_1073;
  reg REGS_1074;
  reg REGS_1075;
  reg REGS_1076;
  reg REGS_1077;
  reg REGS_1078;
  reg REGS_1079;
  reg REGS_1080;
  reg REGS_1081;
  reg REGS_1082;
  reg REGS_1083;
  reg REGS_1084;
  reg REGS_1085;
  reg REGS_1086;
  reg REGS_1087;
  reg REGS_1088;
  reg REGS_1089;
  reg REGS_1090;
  reg REGS_1091;
  reg REGS_1092;
  reg REGS_1093;
  reg REGS_1094;
  reg REGS_1095;
  reg REGS_1096;
  reg REGS_1097;
  reg REGS_1098;
  reg REGS_1099;
  reg REGS_1100;
  reg REGS_1101;
  reg REGS_1102;
  reg REGS_1103;
  reg REGS_1104;
  reg REGS_1105;
  reg REGS_1106;
  reg REGS_1107;
  reg REGS_1108;
  reg REGS_1109;
  reg REGS_1110;
  reg REGS_1111;
  reg REGS_1112;
  reg REGS_1113;
  reg REGS_1114;
  reg REGS_1115;
  reg REGS_1116;
  reg REGS_1117;
  reg REGS_1118;
  reg REGS_1119;
  reg REGS_1120;
  reg REGS_1121;
  reg REGS_1122;
  reg REGS_1123;
  reg REGS_1124;
  reg REGS_1125;
  reg REGS_1126;
  reg REGS_1127;
  reg REGS_1128;
  reg REGS_1129;
  reg REGS_1130;
  reg REGS_1131;
  reg REGS_1132;
  reg REGS_1133;
  reg REGS_1134;
  reg REGS_1135;
  reg REGS_1136;
  reg REGS_1137;
  reg REGS_1138;
  reg REGS_1139;
  reg REGS_1140;
  reg REGS_1141;
  reg REGS_1142;
  reg REGS_1143;
  reg REGS_1144;
  reg REGS_1145;
  reg REGS_1146;
  reg REGS_1147;
  reg REGS_1148;
  reg REGS_1149;
  reg REGS_1150;
  reg REGS_1151;
  reg REGS_1152;
  reg REGS_1153;
  reg REGS_1154;
  reg REGS_1155;
  reg REGS_1156;
  reg REGS_1157;
  reg REGS_1158;
  reg REGS_1159;
  reg REGS_1160;
  reg REGS_1161;
  reg REGS_1162;
  reg REGS_1163;
  reg REGS_1164;
  reg REGS_1165;
  reg REGS_1166;
  reg REGS_1167;
  reg REGS_1168;
  reg REGS_1169;
  reg REGS_1170;
  reg REGS_1171;
  reg REGS_1172;
  reg REGS_1173;
  reg REGS_1174;
  reg REGS_1175;
  reg REGS_1176;
  reg REGS_1177;
  reg REGS_1178;
  reg REGS_1179;
  reg REGS_1180;
  reg REGS_1181;
  reg REGS_1182;
  reg REGS_1183;
  reg REGS_1184;
  reg REGS_1185;
  reg REGS_1186;
  reg REGS_1187;
  reg REGS_1188;
  reg REGS_1189;
  reg REGS_1190;
  reg REGS_1191;
  reg REGS_1192;
  reg REGS_1193;
  reg REGS_1194;
  reg REGS_1195;
  reg REGS_1196;
  reg REGS_1197;
  reg REGS_1198;
  reg REGS_1199;
  reg REGS_1200;
  reg REGS_1201;
  reg REGS_1202;
  reg REGS_1203;
  reg REGS_1204;
  reg REGS_1205;
  reg REGS_1206;
  reg REGS_1207;
  reg REGS_1208;
  reg REGS_1209;
  reg REGS_1210;
  reg REGS_1211;
  reg REGS_1212;
  reg REGS_1213;
  reg REGS_1214;
  reg REGS_1215;
  reg REGS_1216;
  reg REGS_1217;
  reg REGS_1218;
  reg REGS_1219;
  reg REGS_1220;
  reg REGS_1221;
  reg REGS_1222;
  reg REGS_1223;
  reg REGS_1224;
  reg REGS_1225;
  reg REGS_1226;
  reg REGS_1227;
  reg REGS_1228;
  reg REGS_1229;
  reg REGS_1230;
  reg REGS_1231;
  reg REGS_1232;
  reg REGS_1233;
  reg REGS_1234;
  reg REGS_1235;
  reg REGS_1236;
  reg REGS_1237;
  reg REGS_1238;
  reg REGS_1239;
  reg REGS_1240;
  reg REGS_1241;
  reg REGS_1242;
  reg REGS_1243;
  reg REGS_1244;
  reg REGS_1245;
  reg REGS_1246;
  reg REGS_1247;
  reg REGS_1248;
  reg REGS_1249;
  reg REGS_1250;
  reg REGS_1251;
  reg REGS_1252;
  reg REGS_1253;
  reg REGS_1254;
  reg REGS_1255;
  reg REGS_1256;
  reg REGS_1257;
  reg REGS_1258;
  reg REGS_1259;
  reg REGS_1260;
  reg REGS_1261;
  reg REGS_1262;
  reg REGS_1263;
  reg REGS_1264;
  reg REGS_1265;
  reg REGS_1266;
  reg REGS_1267;
  reg REGS_1268;
  reg REGS_1269;
  reg REGS_1270;
  reg REGS_1271;
  reg REGS_1272;
  reg REGS_1273;
  reg REGS_1274;
  reg REGS_1275;
  reg REGS_1276;
  reg REGS_1277;
  reg REGS_1278;
  reg REGS_1279;
  reg REGS_1280;
  reg REGS_1281;
  reg REGS_1282;
  reg REGS_1283;
  reg REGS_1284;
  reg REGS_1285;
  reg REGS_1286;
  reg REGS_1287;
  reg REGS_1288;
  reg REGS_1289;
  reg REGS_1290;
  reg REGS_1291;
  reg REGS_1292;
  reg REGS_1293;
  reg REGS_1294;
  reg REGS_1295;
  reg REGS_1296;
  reg REGS_1297;
  reg REGS_1298;
  reg REGS_1299;
  reg REGS_1300;
  reg REGS_1301;
  reg REGS_1302;
  reg REGS_1303;
  reg REGS_1304;
  reg REGS_1305;
  reg REGS_1306;
  reg REGS_1307;
  reg REGS_1308;
  reg REGS_1309;
  reg REGS_1310;
  reg REGS_1311;
  reg REGS_1312;
  reg REGS_1313;
  reg REGS_1314;
  reg REGS_1315;
  reg REGS_1316;
  reg REGS_1317;
  reg REGS_1318;
  reg REGS_1319;
  reg REGS_1320;
  reg REGS_1321;
  reg REGS_1322;
  reg REGS_1323;
  reg REGS_1324;
  reg REGS_1325;
  reg REGS_1326;
  reg REGS_1327;
  reg REGS_1328;
  reg REGS_1329;
  reg REGS_1330;
  reg REGS_1331;
  reg REGS_1332;
  reg REGS_1333;
  reg REGS_1334;
  reg REGS_1335;
  reg REGS_1336;
  reg REGS_1337;
  reg REGS_1338;
  reg REGS_1339;
  reg REGS_1340;
  reg REGS_1341;
  reg REGS_1342;
  reg REGS_1343;
  reg REGS_1344;
  reg REGS_1345;
  reg REGS_1346;
  reg REGS_1347;
  reg REGS_1348;
  reg REGS_1349;
  reg REGS_1350;
  reg REGS_1351;
  reg REGS_1352;
  reg REGS_1353;
  reg REGS_1354;
  reg REGS_1355;
  reg REGS_1356;
  reg REGS_1357;
  reg REGS_1358;
  reg REGS_1359;
  reg REGS_1360;
  reg REGS_1361;
  reg REGS_1362;
  reg REGS_1363;
  reg REGS_1364;
  reg REGS_1365;
  reg REGS_1366;
  reg REGS_1367;
  reg REGS_1368;
  reg REGS_1369;
  reg REGS_1370;
  reg REGS_1371;
  reg REGS_1372;
  reg REGS_1373;
  reg REGS_1374;
  reg REGS_1375;
  reg REGS_1376;
  reg REGS_1377;
  reg REGS_1378;
  reg REGS_1379;
  reg REGS_1380;
  reg REGS_1381;
  reg REGS_1382;
  reg REGS_1383;
  reg REGS_1384;
  reg REGS_1385;
  reg REGS_1386;
  reg REGS_1387;
  reg REGS_1388;
  reg REGS_1389;
  reg REGS_1390;
  reg REGS_1391;
  reg REGS_1392;
  reg REGS_1393;
  reg REGS_1394;
  reg REGS_1395;
  reg REGS_1396;
  reg REGS_1397;
  reg REGS_1398;
  reg REGS_1399;
  reg REGS_1400;
  reg REGS_1401;
  reg REGS_1402;
  reg REGS_1403;
  reg REGS_1404;
  reg REGS_1405;
  reg REGS_1406;
  reg REGS_1407;
  reg REGS_1408;
  reg REGS_1409;
  reg REGS_1410;
  reg REGS_1411;
  reg REGS_1412;
  reg REGS_1413;
  reg REGS_1414;
  reg REGS_1415;
  reg REGS_1416;
  reg REGS_1417;
  reg REGS_1418;
  reg REGS_1419;
  reg REGS_1420;
  reg REGS_1421;
  reg REGS_1422;
  reg REGS_1423;
  reg REGS_1424;
  reg REGS_1425;
  reg REGS_1426;
  reg REGS_1427;
  reg REGS_1428;
  reg REGS_1429;
  reg REGS_1430;
  reg REGS_1431;
  reg REGS_1432;
  reg REGS_1433;
  reg REGS_1434;
  reg REGS_1435;
  reg REGS_1436;
  reg REGS_1437;
  reg REGS_1438;
  reg REGS_1439;
  reg REGS_1440;
  reg REGS_1441;
  reg REGS_1442;
  reg REGS_1443;
  reg REGS_1444;
  reg REGS_1445;
  reg REGS_1446;
  reg REGS_1447;
  reg REGS_1448;
  reg REGS_1449;
  reg REGS_1450;
  reg REGS_1451;
  reg REGS_1452;
  reg REGS_1453;
  reg REGS_1454;
  reg REGS_1455;
  reg REGS_1456;
  reg REGS_1457;
  reg REGS_1458;
  reg REGS_1459;
  reg REGS_1460;
  reg REGS_1461;
  reg REGS_1462;
  reg REGS_1463;
  reg REGS_1464;
  reg REGS_1465;
  reg REGS_1466;
  reg REGS_1467;
  reg REGS_1468;
  reg REGS_1469;
  reg REGS_1470;
  reg REGS_1471;
  reg REGS_1472;
  reg REGS_1473;
  reg REGS_1474;
  reg REGS_1475;
  reg REGS_1476;
  reg REGS_1477;
  reg REGS_1478;
  reg REGS_1479;
  reg REGS_1480;
  reg REGS_1481;
  reg REGS_1482;
  reg REGS_1483;
  reg REGS_1484;
  reg REGS_1485;
  reg REGS_1486;
  reg REGS_1487;
  reg REGS_1488;
  reg REGS_1489;
  reg REGS_1490;
  reg REGS_1491;
  reg REGS_1492;
  reg REGS_1493;
  reg REGS_1494;
  reg REGS_1495;
  reg REGS_1496;
  reg REGS_1497;
  reg REGS_1498;
  reg REGS_1499;
  reg REGS_1500;
  reg REGS_1501;
  reg REGS_1502;
  reg REGS_1503;
  reg REGS_1504;
  reg REGS_1505;
  reg REGS_1506;
  reg REGS_1507;
  reg REGS_1508;
  reg REGS_1509;
  reg REGS_1510;
  reg REGS_1511;
  reg REGS_1512;
  reg REGS_1513;
  reg REGS_1514;
  reg REGS_1515;
  reg REGS_1516;
  reg REGS_1517;
  reg REGS_1518;
  reg REGS_1519;
  reg REGS_1520;
  reg REGS_1521;
  reg REGS_1522;
  reg REGS_1523;
  reg REGS_1524;
  reg REGS_1525;
  reg REGS_1526;
  reg REGS_1527;
  reg REGS_1528;
  reg REGS_1529;
  reg REGS_1530;
  reg REGS_1531;
  reg REGS_1532;
  reg REGS_1533;
  reg REGS_1534;
  reg REGS_1535;
  reg REGS_1536;
  reg REGS_1537;
  reg REGS_1538;
  reg REGS_1539;
  reg REGS_1540;
  reg REGS_1541;
  reg REGS_1542;
  reg REGS_1543;
  reg REGS_1544;
  reg REGS_1545;
  reg REGS_1546;
  reg REGS_1547;
  reg REGS_1548;
  reg REGS_1549;
  reg REGS_1550;
  reg REGS_1551;
  reg REGS_1552;
  reg REGS_1553;
  reg REGS_1554;
  reg REGS_1555;
  reg REGS_1556;
  reg REGS_1557;
  reg REGS_1558;
  reg REGS_1559;
  reg REGS_1560;
  reg REGS_1561;
  reg REGS_1562;
  reg REGS_1563;
  reg REGS_1564;
  reg REGS_1565;
  reg REGS_1566;
  reg REGS_1567;
  reg REGS_1568;
  reg REGS_1569;
  reg REGS_1570;
  reg REGS_1571;
  reg REGS_1572;
  reg REGS_1573;
  reg REGS_1574;
  reg REGS_1575;
  reg REGS_1576;
  reg REGS_1577;
  reg REGS_1578;
  reg REGS_1579;
  reg REGS_1580;
  reg REGS_1581;
  reg REGS_1582;
  reg REGS_1583;
  reg REGS_1584;
  reg REGS_1585;
  reg REGS_1586;
  reg REGS_1587;
  reg REGS_1588;
  reg REGS_1589;
  reg REGS_1590;
  reg REGS_1591;
  reg REGS_1592;
  reg REGS_1593;
  reg REGS_1594;
  reg REGS_1595;
  reg REGS_1596;
  reg REGS_1597;
  reg REGS_1598;
  reg REGS_1599;
  wire FA_out_0;
  wire FA_out_1;
  wire FA_out_2;
  wire FA_out_3;
  wire FA_out_4;
  wire FA_out_5;
  wire FA_out_6;
  wire FA_out_7;
  wire FA_out_8;
  wire FA_out_9;
  wire FA_out_10;
  wire FA_out_11;
  wire FA_out_12;
  wire FA_out_13;
  wire FA_out_14;
  wire FA_out_15;
  wire FA_out_16;
  wire FA_out_17;
  wire FA_out_18;
  wire FA_out_19;
  wire FA_out_20;
  wire FA_out_21;
  wire FA_out_22;
  wire FA_out_23;
  wire FA_out_24;
  wire FA_out_25;
  wire FA_out_26;
  wire FA_out_27;
  wire FA_out_28;
  wire FA_out_29;
  wire FA_out_30;
  wire FA_out_31;
  wire FA_out_32;
  wire FA_out_33;
  wire FA_out_34;
  wire FA_out_35;
  wire FA_out_36;
  wire FA_out_37;
  wire FA_out_38;
  wire FA_out_39;
  wire FA_out_40;
  wire FA_out_41;
  wire FA_out_42;
  wire FA_out_43;
  wire FA_out_44;
  wire FA_out_45;
  wire FA_out_46;
  wire FA_out_47;
  wire FA_out_48;
  wire FA_out_49;
  wire FA_out_50;
  wire FA_out_51;
  wire FA_out_52;
  wire FA_out_53;
  wire FA_out_54;
  wire FA_out_55;
  wire FA_out_56;
  wire FA_out_57;
  wire FA_out_58;
  wire FA_out_59;
  wire FA_out_60;
  wire FA_out_61;
  wire FA_out_62;
  wire FA_out_63;
  wire FA_out_64;
  wire FA_out_65;
  wire FA_out_66;
  wire FA_out_67;
  wire FA_out_68;
  wire FA_out_69;
  wire FA_out_70;
  wire FA_out_71;
  wire FA_out_72;
  wire FA_out_73;
  wire FA_out_74;
  wire FA_out_75;
  wire FA_out_76;
  wire FA_out_77;
  wire FA_out_78;
  wire FA_out_79;
  wire FA_out_80;
  wire FA_out_81;
  wire FA_out_82;
  wire FA_out_83;
  wire FA_out_84;
  wire FA_out_85;
  wire FA_out_86;
  wire FA_out_87;
  wire FA_out_88;
  wire FA_out_89;
  wire FA_out_90;
  wire FA_out_91;
  wire FA_out_92;
  wire FA_out_93;
  wire FA_out_94;
  wire FA_out_95;
  wire FA_out_96;
  wire FA_out_97;
  wire FA_out_98;
  wire FA_out_99;
  wire FA_out_100;
  wire FA_out_101;
  wire FA_out_102;
  wire FA_out_103;
  wire FA_out_104;
  wire FA_out_105;
  wire FA_out_106;
  wire FA_out_107;
  wire FA_out_108;
  wire FA_out_109;
  wire FA_out_110;
  wire FA_out_111;
  wire FA_out_112;
  wire FA_out_113;
  wire FA_out_114;
  wire FA_out_115;
  wire FA_out_116;
  wire FA_out_117;
  wire FA_out_118;
  wire FA_out_119;
  wire FA_out_120;
  wire FA_out_121;
  wire FA_out_122;
  wire FA_out_123;
  wire FA_out_124;
  wire FA_out_125;
  wire FA_out_126;
  wire FA_out_127;
  wire FA_out_128;
  wire FA_out_129;
  wire FA_out_130;
  wire FA_out_131;
  wire FA_out_132;
  wire FA_out_133;
  wire FA_out_134;
  wire FA_out_135;
  wire FA_out_136;
  wire FA_out_137;
  wire FA_out_138;
  wire FA_out_139;
  wire FA_out_140;
  wire FA_out_141;
  wire FA_out_142;
  wire FA_out_143;
  wire FA_out_144;
  wire FA_out_145;
  wire FA_out_146;
  wire FA_out_147;
  wire FA_out_148;
  wire FA_out_149;
  wire FA_out_150;
  wire FA_out_151;
  wire FA_out_152;
  wire FA_out_153;
  wire FA_out_154;
  wire FA_out_155;
  wire FA_out_156;
  wire FA_out_157;
  wire FA_out_158;
  wire FA_out_159;
  wire FA_out_160;
  wire FA_out_161;
  wire FA_out_162;
  wire FA_out_163;
  wire FA_out_164;
  wire FA_out_165;
  wire FA_out_166;
  wire FA_out_167;
  wire FA_out_168;
  wire FA_out_169;
  wire FA_out_170;
  wire FA_out_171;
  wire FA_out_172;
  wire FA_out_173;
  wire FA_out_174;
  wire FA_out_175;
  wire FA_out_176;
  wire FA_out_177;
  wire FA_out_178;
  wire FA_out_179;
  wire FA_out_180;
  wire FA_out_181;
  wire FA_out_182;
  wire FA_out_183;
  wire FA_out_184;
  wire FA_out_185;
  wire FA_out_186;
  wire FA_out_187;
  wire FA_out_188;
  wire FA_out_189;
  wire FA_out_190;
  wire FA_out_191;
  wire FA_out_192;
  wire FA_out_193;
  wire FA_out_194;
  wire FA_out_195;
  wire FA_out_196;
  wire FA_out_197;
  wire FA_out_198;
  wire FA_out_199;
  wire FA_out_200;
  wire FA_out_201;
  wire FA_out_202;
  wire FA_out_203;
  wire FA_out_204;
  wire FA_out_205;
  wire FA_out_206;
  wire FA_out_207;
  wire FA_out_208;
  wire FA_out_209;
  wire FA_out_210;
  wire FA_out_211;
  wire FA_out_212;
  wire FA_out_213;
  wire FA_out_214;
  wire FA_out_215;
  wire FA_out_216;
  wire FA_out_217;
  wire FA_out_218;
  wire FA_out_219;
  wire FA_out_220;
  wire FA_out_221;
  wire FA_out_222;
  wire FA_out_223;
  wire FA_out_224;
  wire FA_out_225;
  wire FA_out_226;
  wire FA_out_227;
  wire FA_out_228;
  wire FA_out_229;
  wire FA_out_230;
  wire FA_out_231;
  wire FA_out_232;
  wire FA_out_233;
  wire FA_out_234;
  wire FA_out_235;
  wire FA_out_236;
  wire FA_out_237;
  wire FA_out_238;
  wire FA_out_239;
  wire FA_out_240;
  wire FA_out_241;
  wire FA_out_242;
  wire FA_out_243;
  wire FA_out_244;
  wire FA_out_245;
  wire FA_out_246;
  wire FA_out_247;
  wire FA_out_248;
  wire FA_out_249;
  wire FA_out_250;
  wire FA_out_251;
  wire FA_out_252;
  wire FA_out_253;
  wire FA_out_254;
  wire FA_out_255;
  wire FA_out_256;
  wire FA_out_257;
  wire FA_out_258;
  wire FA_out_259;
  wire FA_out_260;
  wire FA_out_261;
  wire FA_out_262;
  wire FA_out_263;
  wire FA_out_264;
  wire FA_out_265;
  wire FA_out_266;
  wire FA_out_267;
  wire FA_out_268;
  wire FA_out_269;
  wire FA_out_270;
  wire FA_out_271;
  wire FA_out_272;
  wire FA_out_273;
  wire FA_out_274;
  wire FA_out_275;
  wire FA_out_276;
  wire FA_out_277;
  wire FA_out_278;
  wire FA_out_279;
  wire FA_out_280;
  wire FA_out_281;
  wire FA_out_282;
  wire FA_out_283;
  wire FA_out_284;
  wire FA_out_285;
  wire FA_out_286;
  wire FA_out_287;
  wire FA_out_288;
  wire FA_out_289;
  wire FA_out_290;
  wire FA_out_291;
  wire FA_out_292;
  wire FA_out_293;
  wire FA_out_294;
  wire FA_out_295;
  wire FA_out_296;
  wire FA_out_297;
  wire FA_out_298;
  wire FA_out_299;
  wire FA_out_300;
  wire FA_out_301;
  wire FA_out_302;
  wire FA_out_303;
  wire FA_out_304;
  wire FA_out_305;
  wire FA_out_306;
  wire FA_out_307;
  wire FA_out_308;
  wire FA_out_309;
  wire FA_out_310;
  wire FA_out_311;
  wire FA_out_312;
  wire FA_out_313;
  wire FA_out_314;
  wire FA_out_315;
  wire FA_out_316;
  wire FA_out_317;
  wire FA_out_318;
  wire FA_out_319;
  wire FA_out_320;
  wire FA_out_321;
  wire FA_out_322;
  wire FA_out_323;
  wire FA_out_324;
  wire FA_out_325;
  wire FA_out_326;
  wire FA_out_327;
  wire FA_out_328;
  wire FA_out_329;
  wire FA_out_330;
  wire FA_out_331;
  wire FA_out_332;
  wire FA_out_333;
  wire FA_out_334;
  wire FA_out_335;
  wire FA_out_336;
  wire FA_out_337;
  wire FA_out_338;
  wire FA_out_339;
  wire FA_out_340;
  wire FA_out_341;
  wire FA_out_342;
  wire FA_out_343;
  wire FA_out_344;
  wire FA_out_345;
  wire FA_out_346;
  wire FA_out_347;
  wire FA_out_348;
  wire FA_out_349;
  wire FA_out_350;
  wire FA_out_351;
  wire FA_out_352;
  wire FA_out_353;
  wire FA_out_354;
  wire FA_out_355;
  wire FA_out_356;
  wire FA_out_357;
  wire FA_out_358;
  wire FA_out_359;
  wire FA_out_360;
  wire FA_out_361;
  wire FA_out_362;
  wire FA_out_363;
  wire FA_out_364;
  wire FA_out_365;
  wire FA_out_366;
  wire FA_out_367;
  wire FA_out_368;
  wire FA_out_369;
  wire FA_out_370;
  wire FA_out_371;
  wire FA_out_372;
  wire FA_out_373;
  wire FA_out_374;
  wire FA_out_375;
  wire FA_out_376;
  wire FA_out_377;
  wire FA_out_378;
  wire FA_out_379;
  wire FA_out_380;
  wire FA_out_381;
  wire FA_out_382;
  wire FA_out_383;
  wire FA_out_384;
  wire FA_out_385;
  wire FA_out_386;
  wire FA_out_387;
  wire FA_out_388;
  wire FA_out_389;
  wire FA_out_390;
  wire FA_out_391;
  wire FA_out_392;
  wire FA_out_393;
  wire FA_out_394;
  wire FA_out_395;
  wire FA_out_396;
  wire FA_out_397;
  wire FA_out_398;
  wire FA_out_399;
  wire FA_out_400;
  wire FA_out_401;
  wire FA_out_402;
  wire FA_out_403;
  wire FA_out_404;
  wire FA_out_405;
  wire FA_out_406;
  wire FA_out_407;
  wire FA_out_408;
  wire FA_out_409;
  wire FA_out_410;
  wire FA_out_411;
  wire FA_out_412;
  wire FA_out_413;
  wire FA_out_414;
  wire FA_out_415;
  wire FA_out_416;
  wire FA_out_417;
  wire FA_out_418;
  wire FA_out_419;
  wire FA_out_420;
  wire FA_out_421;
  wire FA_out_422;
  wire FA_out_423;
  wire FA_out_424;
  wire FA_out_425;
  wire FA_out_426;
  wire FA_out_427;
  wire FA_out_428;
  wire FA_out_429;
  wire FA_out_430;
  wire FA_out_431;
  wire FA_out_432;
  wire FA_out_433;
  wire FA_out_434;
  wire FA_out_435;
  wire FA_out_436;
  wire FA_out_437;
  wire FA_out_438;
  wire FA_out_439;
  wire FA_out_440;
  wire FA_out_441;
  wire FA_out_442;
  wire FA_out_443;
  wire FA_out_444;
  wire FA_out_445;
  wire FA_out_446;
  wire FA_out_447;
  wire FA_out_448;
  wire FA_out_449;
  wire FA_out_450;
  wire FA_out_451;
  wire FA_out_452;
  wire FA_out_453;
  wire FA_out_454;
  wire FA_out_455;
  wire FA_out_456;
  wire FA_out_457;
  wire FA_out_458;
  wire FA_out_459;
  wire FA_out_460;
  wire FA_out_461;
  wire FA_out_462;
  wire FA_out_463;
  wire FA_out_464;
  wire FA_out_465;
  wire FA_out_466;
  wire FA_out_467;
  wire FA_out_468;
  wire FA_out_469;
  wire FA_out_470;
  wire FA_out_471;
  wire FA_out_472;
  wire FA_out_473;
  wire FA_out_474;
  wire FA_out_475;
  wire FA_out_476;
  wire FA_out_477;
  wire FA_out_478;
  wire FA_out_479;
  wire FA_out_480;
  wire FA_out_481;
  wire FA_out_482;
  wire FA_out_483;
  wire FA_out_484;
  wire FA_out_485;
  wire FA_out_486;
  wire FA_out_487;
  wire FA_out_488;
  wire FA_out_489;
  wire FA_out_490;
  wire FA_out_491;
  wire FA_out_492;
  wire FA_out_493;
  wire FA_out_494;
  wire FA_out_495;
  wire FA_out_496;
  wire FA_out_497;
  wire FA_out_498;
  wire FA_out_499;
  wire FA_out_500;
  wire FA_out_501;
  wire FA_out_502;
  wire FA_out_503;
  wire FA_out_504;
  wire FA_out_505;
  wire FA_out_506;
  wire FA_out_507;
  wire FA_out_508;
  wire FA_out_509;
  wire FA_out_510;
  wire FA_out_511;
  wire FA_out_512;
  wire FA_out_513;
  wire FA_out_514;
  wire FA_out_515;
  wire FA_out_516;
  wire FA_out_517;
  wire FA_out_518;
  wire FA_out_519;
  wire FA_out_520;
  wire FA_out_521;
  wire FA_out_522;
  wire FA_out_523;
  wire FA_out_524;
  wire FA_out_525;
  wire FA_out_526;
  wire FA_out_527;
  wire FA_out_528;
  wire FA_out_529;
  wire FA_out_530;
  wire FA_out_531;
  wire FA_out_532;
  wire FA_out_533;
  wire FA_out_534;
  wire FA_out_535;
  wire FA_out_536;
  wire FA_out_537;
  wire FA_out_538;
  wire FA_out_539;
  wire FA_out_540;
  wire FA_out_541;
  wire FA_out_542;
  wire FA_out_543;
  wire FA_out_544;
  wire FA_out_545;
  wire FA_out_546;
  wire FA_out_547;
  wire FA_out_548;
  wire FA_out_549;
  wire FA_out_550;
  wire FA_out_551;
  wire FA_out_552;
  wire FA_out_553;
  wire FA_out_554;
  wire FA_out_555;
  wire FA_out_556;
  wire FA_out_557;
  wire FA_out_558;
  wire FA_out_559;
  wire FA_out_560;
  wire FA_out_561;
  wire FA_out_562;
  wire FA_out_563;
  wire FA_out_564;
  wire FA_out_565;
  wire FA_out_566;
  wire FA_out_567;
  wire FA_out_568;
  wire FA_out_569;
  wire FA_out_570;
  wire FA_out_571;
  wire FA_out_572;
  wire FA_out_573;
  wire FA_out_574;
  wire FA_out_575;
  wire FA_out_576;
  wire FA_out_577;
  wire FA_out_578;
  wire FA_out_579;
  wire FA_out_580;
  wire FA_out_581;
  wire FA_out_582;
  wire FA_out_583;
  wire FA_out_584;
  wire FA_out_585;
  wire FA_out_586;
  wire FA_out_587;
  wire FA_out_588;
  wire FA_out_589;
  wire FA_out_590;
  wire FA_out_591;
  wire FA_out_592;
  wire FA_out_593;
  wire FA_out_594;
  wire FA_out_595;
  wire FA_out_596;
  wire FA_out_597;
  wire FA_out_598;
  wire FA_out_599;
  wire FA_out_600;
  wire FA_out_601;
  wire FA_out_602;
  wire FA_out_603;
  wire FA_out_604;
  wire FA_out_605;
  wire FA_out_606;
  wire FA_out_607;
  wire FA_out_608;
  wire FA_out_609;
  wire FA_out_610;
  wire FA_out_611;
  wire FA_out_612;
  wire FA_out_613;
  wire FA_out_614;
  wire FA_out_615;
  wire FA_out_616;
  wire FA_out_617;
  wire FA_out_618;
  wire FA_out_619;
  wire FA_out_620;
  wire FA_out_621;
  wire FA_out_622;
  wire FA_out_623;
  wire FA_out_624;
  wire FA_out_625;
  wire FA_out_626;
  wire FA_out_627;
  wire FA_out_628;
  wire FA_out_629;
  wire FA_out_630;
  wire FA_out_631;
  wire FA_out_632;
  wire FA_out_633;
  wire FA_out_634;
  wire FA_out_635;
  wire FA_out_636;
  wire FA_out_637;
  wire FA_out_638;
  wire FA_out_639;
  wire FA_out_640;
  wire FA_out_641;
  wire FA_out_642;
  wire FA_out_643;
  wire FA_out_644;
  wire FA_out_645;
  wire FA_out_646;
  wire FA_out_647;
  wire FA_out_648;
  wire FA_out_649;
  wire FA_out_650;
  wire FA_out_651;
  wire FA_out_652;
  wire FA_out_653;
  wire FA_out_654;
  wire FA_out_655;
  wire FA_out_656;
  wire FA_out_657;
  wire FA_out_658;
  wire FA_out_659;
  wire FA_out_660;
  wire FA_out_661;
  wire FA_out_662;
  wire FA_out_663;
  wire FA_out_664;
  wire FA_out_665;
  wire FA_out_666;
  wire FA_out_667;
  wire FA_out_668;
  wire FA_out_669;
  wire FA_out_670;
  wire FA_out_671;
  wire FA_out_672;
  wire FA_out_673;
  wire FA_out_674;
  wire FA_out_675;
  wire FA_out_676;
  wire FA_out_677;
  wire FA_out_678;
  wire FA_out_679;
  wire FA_out_680;
  wire FA_out_681;
  wire FA_out_682;
  wire FA_out_683;
  wire FA_out_684;
  wire FA_out_685;
  wire FA_out_686;
  wire FA_out_687;
  wire FA_out_688;
  wire FA_out_689;
  wire FA_out_690;
  wire FA_out_691;
  wire FA_out_692;
  wire FA_out_693;
  wire FA_out_694;
  wire FA_out_695;
  wire FA_out_696;
  wire FA_out_697;
  wire FA_out_698;
  wire FA_out_699;
  wire FA_out_700;
  wire FA_out_701;
  wire FA_out_702;
  wire FA_out_703;
  wire FA_out_704;
  wire FA_out_705;
  wire FA_out_706;
  wire FA_out_707;
  wire FA_out_708;
  wire FA_out_709;
  wire FA_out_710;
  wire FA_out_711;
  wire FA_out_712;
  wire FA_out_713;
  wire FA_out_714;
  wire FA_out_715;
  wire FA_out_716;
  wire FA_out_717;
  wire FA_out_718;
  wire FA_out_719;
  wire FA_out_720;
  wire FA_out_721;
  wire FA_out_722;
  wire FA_out_723;
  wire FA_out_724;
  wire FA_out_725;
  wire FA_out_726;
  wire FA_out_727;
  wire FA_out_728;
  wire FA_out_729;
  wire FA_out_730;
  wire FA_out_731;
  wire FA_out_732;
  wire FA_out_733;
  wire FA_out_734;
  wire FA_out_735;
  wire FA_out_736;
  wire FA_out_737;
  wire FA_out_738;
  wire FA_out_739;
  wire FA_out_740;
  wire FA_out_741;
  wire FA_out_742;
  wire FA_out_743;
  wire FA_out_744;
  wire FA_out_745;
  wire FA_out_746;
  wire FA_out_747;
  wire FA_out_748;
  wire FA_out_749;
  wire FA_out_750;
  wire FA_out_751;
  wire FA_out_752;
  wire FA_out_753;
  wire FA_out_754;
  wire FA_out_755;
  wire FA_out_756;
  wire FA_out_757;
  wire FA_out_758;
  wire FA_out_759;
  wire FA_out_760;
  wire FA_out_761;
  wire FA_out_762;
  wire FA_out_763;
  wire FA_out_764;
  wire FA_out_765;
  wire FA_out_766;
  wire FA_out_767;
  wire FA_out_768;
  wire FA_out_769;
  wire FA_out_770;
  wire FA_out_771;
  wire FA_out_772;
  wire FA_out_773;
  wire FA_out_774;
  wire FA_out_775;
  wire FA_out_776;
  wire FA_out_777;
  wire FA_out_778;
  wire FA_out_779;
  wire FA_out_780;
  wire FA_out_781;
  wire FA_out_782;
  wire FA_out_783;
  wire FA_out_784;
  wire FA_out_785;
  wire FA_out_786;
  wire FA_out_787;
  wire FA_out_788;
  wire FA_out_789;
  wire FA_out_790;
  wire FA_out_791;
  wire FA_out_792;
  wire FA_out_793;
  wire FA_out_794;
  wire FA_out_795;
  wire FA_out_796;
  wire FA_out_797;
  wire FA_out_798;
  wire FA_out_799;
  wire FA_out_800;
  wire FA_out_801;
  wire FA_out_802;
  wire FA_out_803;
  wire FA_out_804;
  wire FA_out_805;
  wire FA_out_806;
  wire FA_out_807;
  wire FA_out_808;
  wire FA_out_809;
  wire FA_out_810;
  wire FA_out_811;
  wire FA_out_812;
  wire FA_out_813;
  wire FA_out_814;
  wire FA_out_815;
  wire FA_out_816;
  wire FA_out_817;
  wire FA_out_818;
  wire FA_out_819;
  wire FA_out_820;
  wire FA_out_821;
  wire FA_out_822;
  wire FA_out_823;
  wire FA_out_824;
  wire FA_out_825;
  wire FA_out_826;
  wire FA_out_827;
  wire FA_out_828;
  wire FA_out_829;
  wire FA_out_830;
  wire FA_out_831;
  wire FA_out_832;
  wire FA_out_833;
  wire FA_out_834;
  wire FA_out_835;
  wire FA_out_836;
  wire FA_out_837;
  wire FA_out_838;
  wire FA_out_839;
  wire FA_out_840;
  wire FA_out_841;
  wire FA_out_842;
  wire FA_out_843;
  wire FA_out_844;
  wire FA_out_845;
  wire FA_out_846;
  wire FA_out_847;
  wire FA_out_848;
  wire FA_out_849;
  wire FA_out_850;
  wire FA_out_851;
  wire FA_out_852;
  wire FA_out_853;
  wire FA_out_854;
  wire FA_out_855;
  wire FA_out_856;
  wire FA_out_857;
  wire FA_out_858;
  wire FA_out_859;
  wire FA_out_860;
  wire FA_out_861;
  wire FA_out_862;
  wire FA_out_863;
  wire FA_out_864;
  wire FA_out_865;
  wire FA_out_866;
  wire FA_out_867;
  wire FA_out_868;
  wire FA_out_869;
  wire FA_out_870;
  wire FA_out_871;
  wire FA_out_872;
  wire FA_out_873;
  wire FA_out_874;
  wire FA_out_875;
  wire FA_out_876;
  wire FA_out_877;
  wire FA_out_878;
  wire FA_out_879;
  wire FA_out_880;
  wire FA_out_881;
  wire FA_out_882;
  wire FA_out_883;
  wire FA_out_884;
  wire FA_out_885;
  wire FA_out_886;
  wire FA_out_887;
  wire FA_out_888;
  wire FA_out_889;
  wire FA_out_890;
  wire FA_out_891;
  wire FA_out_892;
  wire FA_out_893;
  wire FA_out_894;
  wire FA_out_895;
  wire FA_out_896;
  wire FA_out_897;
  wire FA_out_898;
  wire FA_out_899;
  wire FA_out_900;
  wire FA_out_901;
  wire FA_out_902;
  wire FA_out_903;
  wire FA_out_904;
  wire FA_out_905;
  wire FA_out_906;
  wire FA_out_907;
  wire FA_out_908;
  wire FA_out_909;
  wire FA_out_910;
  wire FA_out_911;
  wire FA_out_912;
  wire FA_out_913;
  wire FA_out_914;
  wire FA_out_915;
  wire FA_out_916;
  wire FA_out_917;
  wire FA_out_918;
  wire FA_out_919;
  wire FA_out_920;
  wire FA_out_921;
  wire FA_out_922;
  wire FA_out_923;
  wire FA_out_924;
  wire FA_out_925;
  wire FA_out_926;
  wire FA_out_927;
  wire FA_out_928;
  wire FA_out_929;
  wire FA_out_930;
  wire FA_out_931;
  wire FA_out_932;
  wire FA_out_933;
  wire FA_out_934;
  wire FA_out_935;
  wire FA_out_936;
  wire FA_out_937;
  wire FA_out_938;
  wire FA_out_939;
  wire FA_out_940;
  wire FA_out_941;
  wire FA_out_942;
  wire FA_out_943;
  wire FA_out_944;
  wire FA_out_945;
  wire FA_out_946;
  wire FA_out_947;
  wire FA_out_948;
  wire FA_out_949;
  wire FA_out_950;
  wire FA_out_951;
  wire FA_out_952;
  wire FA_out_953;
  wire FA_out_954;
  wire FA_out_955;
  wire FA_out_956;
  wire FA_out_957;
  wire FA_out_958;
  wire FA_out_959;
  wire FA_out_960;
  wire FA_out_961;
  wire FA_out_962;
  wire FA_out_963;
  wire FA_out_964;
  wire FA_out_965;
  wire FA_out_966;
  wire FA_out_967;
  wire FA_out_968;
  wire FA_out_969;
  wire FA_out_970;
  wire FA_out_971;
  wire FA_out_972;
  wire FA_out_973;
  wire FA_out_974;
  wire FA_out_975;
  wire FA_out_976;
  wire FA_out_977;
  wire FA_out_978;
  wire FA_out_979;
  wire FA_out_980;
  wire FA_out_981;
  wire FA_out_982;
  wire FA_out_983;
  wire FA_out_984;
  wire FA_out_985;
  wire FA_out_986;
  wire FA_out_987;
  wire FA_out_988;
  wire FA_out_989;
  wire FA_out_990;
  wire FA_out_991;
  wire FA_out_992;
  wire FA_out_993;
  wire FA_out_994;
  wire FA_out_995;
  wire FA_out_996;
  wire FA_out_997;
  wire FA_out_998;
  wire FA_out_999;
  wire FA_out_1000;
  wire FA_out_1001;
  wire FA_out_1002;
  wire FA_out_1003;
  wire FA_out_1004;
  wire FA_out_1005;
  wire FA_out_1006;
  wire FA_out_1007;
  wire FA_out_1008;
  wire FA_out_1009;
  wire FA_out_1010;
  wire FA_out_1011;
  wire FA_out_1012;
  wire FA_out_1013;
  wire FA_out_1014;
  wire FA_out_1015;
  wire FA_out_1016;
  wire FA_out_1017;
  wire FA_out_1018;
  wire FA_out_1019;
  wire FA_out_1020;
  wire FA_out_1021;
  wire FA_out_1022;
  wire FA_out_1023;
  wire FA_out_1024;
  wire FA_out_1025;
  wire FA_out_1026;
  wire FA_out_1027;
  wire FA_out_1028;
  wire FA_out_1029;
  wire FA_out_1030;
  wire FA_out_1031;
  wire FA_out_1032;
  wire FA_out_1033;
  wire FA_out_1034;
  wire FA_out_1035;
  wire FA_out_1036;
  wire FA_out_1037;
  wire FA_out_1038;
  wire FA_out_1039;
  wire FA_out_1040;
  wire FA_out_1041;
  wire FA_out_1042;
  wire FA_out_1043;
  wire FA_out_1044;
  wire FA_out_1045;
  wire FA_out_1046;
  wire FA_out_1047;
  wire FA_out_1048;
  wire FA_out_1049;
  wire FA_out_1050;
  wire FA_out_1051;
  wire FA_out_1052;
  wire FA_out_1053;
  wire FA_out_1054;
  wire FA_out_1055;
  wire FA_out_1056;
  wire FA_out_1057;
  wire FA_out_1058;
  wire FA_out_1059;
  wire FA_out_1060;
  wire FA_out_1061;
  wire FA_out_1062;
  wire FA_out_1063;
  wire FA_out_1064;
  wire FA_out_1065;
  wire FA_out_1066;
  wire FA_out_1067;
  wire FA_out_1068;
  wire FA_out_1069;
  wire FA_out_1070;
  wire FA_out_1071;
  wire FA_out_1072;
  wire FA_out_1073;
  wire FA_out_1074;
  wire FA_out_1075;
  wire FA_out_1076;
  wire FA_out_1077;
  wire FA_out_1078;
  wire FA_out_1079;
  wire FA_out_1080;
  wire FA_out_1081;
  wire FA_out_1082;
  wire FA_out_1083;
  wire FA_out_1084;
  wire FA_out_1085;
  wire FA_out_1086;
  wire FA_out_1087;
  wire FA_out_1088;
  wire FA_out_1089;
  wire FA_out_1090;
  wire FA_out_1091;
  wire FA_out_1092;
  wire FA_out_1093;
  wire FA_out_1094;
  wire FA_out_1095;
  wire FA_out_1096;
  wire FA_out_1097;
  wire FA_out_1098;
  wire FA_out_1099;
  wire FA_out_1100;
  wire FA_out_1101;
  wire FA_out_1102;
  wire FA_out_1103;
  wire FA_out_1104;
  wire FA_out_1105;
  wire FA_out_1106;
  wire FA_out_1107;
  wire FA_out_1108;
  wire FA_out_1109;
  wire FA_out_1110;
  wire FA_out_1111;
  wire FA_out_1112;
  wire FA_out_1113;
  wire FA_out_1114;
  wire FA_out_1115;
  wire FA_out_1116;
  wire FA_out_1117;
  wire FA_out_1118;
  wire FA_out_1119;
  wire FA_out_1120;
  wire FA_out_1121;
  wire FA_out_1122;
  wire FA_out_1123;
  wire FA_out_1124;
  wire FA_out_1125;
  wire FA_out_1126;
  wire FA_out_1127;
  wire FA_out_1128;
  wire FA_out_1129;
  wire FA_out_1130;
  wire FA_out_1131;
  wire FA_out_1132;
  wire FA_out_1133;
  wire FA_out_1134;
  wire FA_out_1135;
  wire FA_out_1136;
  wire FA_out_1137;
  wire FA_out_1138;
  wire FA_out_1139;
  wire FA_out_1140;
  wire FA_out_1141;
  wire FA_out_1142;
  wire FA_out_1143;
  wire FA_out_1144;
  wire FA_out_1145;
  wire FA_out_1146;
  wire FA_out_1147;
  wire FA_out_1148;
  wire FA_out_1149;
  wire FA_out_1150;
  wire FA_out_1151;
  wire FA_out_1152;
  wire FA_out_1153;
  wire FA_out_1154;
  wire FA_out_1155;
  wire FA_out_1156;
  wire FA_out_1157;
  wire FA_out_1158;
  wire FA_out_1159;
  wire FA_out_1160;
  wire FA_out_1161;
  wire FA_out_1162;
  wire FA_out_1163;
  wire FA_out_1164;
  wire FA_out_1165;
  wire FA_out_1166;
  wire FA_out_1167;
  wire FA_out_1168;
  wire FA_out_1169;
  wire FA_out_1170;
  wire FA_out_1171;
  wire FA_out_1172;
  wire FA_out_1173;
  wire FA_out_1174;
  wire FA_out_1175;
  wire FA_out_1176;
  wire FA_out_1177;
  wire FA_out_1178;
  wire FA_out_1179;
  wire FA_out_1180;
  wire FA_out_1181;
  wire FA_out_1182;
  wire FA_out_1183;
  wire FA_out_1184;
  wire FA_out_1185;
  wire FA_out_1186;
  wire FA_out_1187;
  wire FA_out_1188;
  wire FA_out_1189;
  wire FA_out_1190;
  wire FA_out_1191;
  wire FA_out_1192;
  wire FA_out_1193;
  wire FA_out_1194;
  wire FA_out_1195;
  wire FA_out_1196;
  wire FA_out_1197;
  wire FA_out_1198;
  wire FA_out_1199;
  wire FA_out_1200;
  wire FA_out_1201;
  wire FA_out_1202;
  wire FA_out_1203;
  wire FA_out_1204;
  wire FA_out_1205;
  wire FA_out_1206;
  wire FA_out_1207;
  wire FA_out_1208;
  wire FA_out_1209;
  wire FA_out_1210;
  wire FA_out_1211;
  wire FA_out_1212;
  wire FA_out_1213;
  wire FA_out_1214;
  wire FA_out_1215;
  wire FA_out_1216;
  wire FA_out_1217;
  wire FA_out_1218;
  wire FA_out_1219;
  wire FA_out_1220;
  wire FA_out_1221;
  wire FA_out_1222;
  wire FA_out_1223;
  wire FA_out_1224;
  wire FA_out_1225;
  wire FA_out_1226;
  wire FA_out_1227;
  wire FA_out_1228;
  wire FA_out_1229;
  wire FA_out_1230;
  wire FA_out_1231;
  wire FA_out_1232;
  wire FA_out_1233;
  wire FA_out_1234;
  wire FA_out_1235;
  wire FA_out_1236;
  wire FA_out_1237;
  wire FA_out_1238;
  wire FA_out_1239;
  wire FA_out_1240;
  wire FA_out_1241;
  wire FA_out_1242;
  wire FA_out_1243;
  wire FA_out_1244;
  wire FA_out_1245;
  wire FA_out_1246;
  wire FA_out_1247;
  wire FA_out_1248;
  wire FA_out_1249;
  wire FA_out_1250;
  wire FA_out_1251;
  wire FA_out_1252;
  wire FA_out_1253;
  wire FA_out_1254;
  wire FA_out_1255;
  wire FA_out_1256;
  wire FA_out_1257;
  wire FA_out_1258;
  wire FA_out_1259;
  wire FA_out_1260;
  wire FA_out_1261;
  wire FA_out_1262;
  wire FA_out_1263;
  wire FA_out_1264;
  wire FA_out_1265;
  wire FA_out_1266;
  wire FA_out_1267;
  wire FA_out_1268;
  wire FA_out_1269;
  wire FA_out_1270;
  wire FA_out_1271;
  wire FA_out_1272;
  wire FA_out_1273;
  wire FA_out_1274;
  wire FA_out_1275;
  wire FA_out_1276;
  wire FA_out_1277;
  wire FA_out_1278;
  wire FA_out_1279;
  wire FA_out_1280;
  wire FA_out_1281;
  wire FA_out_1282;
  wire FA_out_1283;
  wire FA_out_1284;
  wire FA_out_1285;
  wire FA_out_1286;
  wire FA_out_1287;
  wire FA_out_1288;
  wire FA_out_1289;
  wire FA_out_1290;
  wire FA_out_1291;
  wire FA_out_1292;
  wire FA_out_1293;
  wire FA_out_1294;
  wire FA_out_1295;
  wire FA_out_1296;
  wire FA_out_1297;
  wire FA_out_1298;
  wire FA_out_1299;
  wire FA_out_1300;
  wire FA_out_1301;
  wire FA_out_1302;
  wire FA_out_1303;
  wire FA_out_1304;
  wire FA_out_1305;
  wire FA_out_1306;
  wire FA_out_1307;
  wire FA_out_1308;
  wire FA_out_1309;
  wire FA_out_1310;
  wire FA_out_1311;
  wire FA_out_1312;
  wire FA_out_1313;
  wire FA_out_1314;
  wire FA_out_1315;
  wire FA_out_1316;
  wire FA_out_1317;
  wire FA_out_1318;
  wire FA_out_1319;
  wire FA_out_1320;
  wire FA_out_1321;
  wire FA_out_1322;
  wire FA_out_1323;
  wire FA_out_1324;
  wire FA_out_1325;
  wire FA_out_1326;
  wire FA_out_1327;
  wire FA_out_1328;
  wire FA_out_1329;
  wire FA_out_1330;
  wire FA_out_1331;
  wire FA_out_1332;
  wire FA_out_1333;
  wire FA_out_1334;
  wire FA_out_1335;
  wire FA_out_1336;
  wire FA_out_1337;
  wire FA_out_1338;
  wire FA_out_1339;
  wire FA_out_1340;
  wire FA_out_1341;
  wire FA_out_1342;
  wire FA_out_1343;
  wire FA_out_1344;
  wire FA_out_1345;
  wire FA_out_1346;
  wire FA_out_1347;
  wire FA_out_1348;
  wire FA_out_1349;
  wire FA_out_1350;
  wire FA_out_1351;
  wire FA_out_1352;
  wire FA_out_1353;
  wire FA_out_1354;
  wire FA_out_1355;
  wire FA_out_1356;
  wire FA_out_1357;
  wire FA_out_1358;
  wire FA_out_1359;
  wire FA_out_1360;
  wire FA_out_1361;
  wire FA_out_1362;
  wire FA_out_1363;
  wire FA_out_1364;
  wire FA_out_1365;
  wire FA_out_1366;
  wire FA_out_1367;
  wire FA_out_1368;
  wire FA_out_1369;
  wire FA_out_1370;
  wire FA_out_1371;
  wire FA_out_1372;
  wire FA_out_1373;
  wire FA_out_1374;
  wire FA_out_1375;
  wire FA_out_1376;
  wire FA_out_1377;
  wire FA_out_1378;
  wire FA_out_1379;
  wire FA_out_1380;
  wire FA_out_1381;
  wire FA_out_1382;
  wire FA_out_1383;
  wire FA_out_1384;
  wire FA_out_1385;
  wire FA_out_1386;
  wire FA_out_1387;
  wire FA_out_1388;
  wire FA_out_1389;
  wire FA_out_1390;
  wire FA_out_1391;
  wire FA_out_1392;
  wire FA_out_1393;
  wire FA_out_1394;
  wire FA_out_1395;
  wire FA_out_1396;
  wire FA_out_1397;
  wire FA_out_1398;
  wire FA_out_1399;
  wire FA_out_1400;
  wire FA_out_1401;
  wire FA_out_1402;
  wire FA_out_1403;
  wire FA_out_1404;
  wire FA_out_1405;
  wire FA_out_1406;
  wire FA_out_1407;
  wire FA_out_1408;
  wire FA_out_1409;
  wire FA_out_1410;
  wire FA_out_1411;
  wire FA_out_1412;
  wire FA_out_1413;
  wire FA_out_1414;
  wire FA_out_1415;
  wire FA_out_1416;
  wire FA_out_1417;
  wire FA_out_1418;
  wire FA_out_1419;
  wire FA_out_1420;
  wire FA_out_1421;
  wire FA_out_1422;
  wire FA_out_1423;
  wire FA_out_1424;
  wire FA_out_1425;
  wire FA_out_1426;
  wire FA_out_1427;
  wire FA_out_1428;
  wire FA_out_1429;
  wire FA_out_1430;
  wire FA_out_1431;
  wire FA_out_1432;
  wire FA_out_1433;
  wire FA_out_1434;
  wire FA_out_1435;
  wire FA_out_1436;
  wire FA_out_1437;
  wire FA_out_1438;
  wire FA_out_1439;
  wire FA_out_1440;
  wire FA_out_1441;
  wire FA_out_1442;
  wire FA_out_1443;
  wire FA_out_1444;
  wire FA_out_1445;
  wire FA_out_1446;
  wire FA_out_1447;
  wire FA_out_1448;
  wire FA_out_1449;
  wire FA_out_1450;
  wire FA_out_1451;
  wire FA_out_1452;
  wire FA_out_1453;
  wire FA_out_1454;
  wire FA_out_1455;
  wire FA_out_1456;
  wire FA_out_1457;
  wire FA_out_1458;
  wire FA_out_1459;
  wire FA_out_1460;
  wire FA_out_1461;
  wire FA_out_1462;
  wire FA_out_1463;
  wire FA_out_1464;
  wire FA_out_1465;
  wire FA_out_1466;
  wire FA_out_1467;
  wire FA_out_1468;
  wire FA_out_1469;
  wire FA_out_1470;
  wire FA_out_1471;
  wire FA_out_1472;
  wire FA_out_1473;
  wire FA_out_1474;
  wire FA_out_1475;
  wire FA_out_1476;
  wire FA_out_1477;
  wire FA_out_1478;
  wire FA_out_1479;
  wire FA_out_1480;
  wire FA_out_1481;
  wire FA_out_1482;
  wire FA_out_1483;
  wire FA_out_1484;
  wire FA_out_1485;
  wire FA_out_1486;
  wire FA_out_1487;
  wire FA_out_1488;
  wire FA_out_1489;
  wire FA_out_1490;
  wire FA_out_1491;
  wire FA_out_1492;
  wire FA_out_1493;
  wire FA_out_1494;
  wire FA_out_1495;
  wire FA_out_1496;
  wire FA_out_1497;
  wire FA_out_1498;
  wire FA_out_1499;
  wire FA_out_1500;
  wire FA_out_1501;
  wire FA_out_1502;
  wire FA_out_1503;
  wire FA_out_1504;
  wire FA_out_1505;
  wire FA_out_1506;
  wire FA_out_1507;
  wire FA_out_1508;
  wire FA_out_1509;
  wire FA_out_1510;
  wire FA_out_1511;
  wire FA_out_1512;
  wire FA_out_1513;
  wire FA_out_1514;
  wire FA_out_1515;
  wire FA_out_1516;
  wire FA_out_1517;
  wire FA_out_1518;
  wire FA_out_1519;
  wire FA_out_1520;
  wire FA_out_1521;
  wire FA_out_1522;
  wire FA_out_1523;
  wire FA_out_1524;
  wire FA_out_1525;
  wire FA_out_1526;
  wire FA_out_1527;
  wire FA_out_1528;
  wire FA_out_1529;
  wire FA_out_1530;
  wire FA_out_1531;
  wire FA_out_1532;
  wire FA_out_1533;
  wire FA_out_1534;
  wire FA_out_1535;
  wire FA_out_1536;
  wire FA_out_1537;
  wire FA_out_1538;
  wire FA_out_1539;
  wire FA_out_1540;
  wire FA_out_1541;
  wire FA_out_1542;
  wire FA_out_1543;
  wire FA_out_1544;
  wire FA_out_1545;
  wire FA_out_1546;
  wire FA_out_1547;
  wire FA_out_1548;
  wire FA_out_1549;
  wire FA_out_1550;
  wire FA_out_1551;
  wire FA_out_1552;
  wire FA_out_1553;
  wire FA_out_1554;
  wire FA_out_1555;
  wire FA_out_1556;
  wire FA_out_1557;
  wire FA_out_1558;
  wire FA_out_1559;
  wire FA_out_1560;
  wire FA_out_1561;
  wire FA_out_1562;
  wire FA_out_1563;
  wire FA_out_1564;
  wire FA_out_1565;
  wire FA_out_1566;
  wire FA_out_1567;
  wire FA_out_1568;
  wire FA_out_1569;
  wire FA_out_1570;
  wire FA_out_1571;
  wire FA_out_1572;
  wire FA_out_1573;
  wire FA_out_1574;
  wire FA_out_1575;
  wire FA_out_1576;
  wire FA_out_1577;
  wire FA_out_1578;
  wire FA_out_1579;
  wire FA_out_1580;
  wire FA_out_1581;
  wire FA_out_1582;
  wire FA_out_1583;
  wire FA_out_1584;
  wire FA_out_1585;
  wire FA_out_1586;
  wire FA_out_1587;
  wire FA_out_1588;
  wire FA_out_1589;
  wire FA_out_1590;
  wire FA_out_1591;
  wire FA_out_1592;
  wire FA_out_1593;
  wire FA_out_1594;
  wire FA_out_1595;
  wire FA_out_1596;
  wire FA_out_1597;
  wire FA_out_1598;
  wire FA_out_1599;
  wire FA_out_1600;
  wire FA_out_1601;
  wire FA_out_1602;
  wire FA_out_1603;
  wire FA_out_1604;
  wire FA_out_1605;
  wire FA_out_1606;
  wire FA_out_1607;
  wire FA_out_1608;
  wire FA_out_1609;
  wire FA_out_1610;
  wire FA_out_1611;
  wire FA_out_1612;
  wire FA_out_1613;
  wire FA_out_1614;
  wire FA_out_1615;
  wire FA_out_1616;
  wire FA_out_1617;
  wire FA_out_1618;
  wire FA_out_1619;
  wire FA_out_1620;
  wire FA_out_1621;
  wire FA_out_1622;
  wire FA_out_1623;
  wire FA_out_1624;
  wire FA_out_1625;
  wire FA_out_1626;
  wire FA_out_1627;
  wire FA_out_1628;
  wire FA_out_1629;
  wire FA_out_1630;
  wire FA_out_1631;
  wire FA_out_1632;
  wire FA_out_1633;
  wire FA_out_1634;
  wire FA_out_1635;
  wire FA_out_1636;
  wire FA_out_1637;
  wire FA_out_1638;
  wire FA_out_1639;
  wire FA_out_1640;
  wire FA_out_1641;
  wire FA_out_1642;
  wire FA_out_1643;
  wire FA_out_1644;
  wire FA_out_1645;
  wire FA_out_1646;
  wire FA_out_1647;
  wire FA_out_1648;
  wire FA_out_1649;
  wire FA_out_1650;
  wire FA_out_1651;
  wire FA_out_1652;
  wire FA_out_1653;
  wire FA_out_1654;
  wire FA_out_1655;
  wire FA_out_1656;
  wire FA_out_1657;
  wire FA_out_1658;
  wire FA_out_1659;
  wire FA_out_1660;
  wire FA_out_1661;
  wire FA_out_1662;
  wire FA_out_1663;
  wire FA_out_1664;
  wire FA_out_1665;
  wire FA_out_1666;
  wire FA_out_1667;
  wire FA_out_1668;
  wire FA_out_1669;
  wire FA_out_1670;
  wire FA_out_1671;
  wire FA_out_1672;
  wire FA_out_1673;
  wire FA_out_1674;
  wire FA_out_1675;
  wire FA_out_1676;
  wire FA_out_1677;
  wire FA_out_1678;
  wire FA_out_1679;
  wire FA_out_1680;
  wire FA_out_1681;
  wire FA_out_1682;
  wire FA_out_1683;
  wire FA_out_1684;
  wire FA_out_1685;
  wire FA_out_1686;
  wire FA_out_1687;
  wire FA_out_1688;
  wire FA_out_1689;
  wire FA_out_1690;
  wire FA_out_1691;
  wire FA_out_1692;
  wire FA_out_1693;
  wire FA_out_1694;
  wire FA_out_1695;
  wire FA_out_1696;
  wire FA_out_1697;
  wire FA_out_1698;
  wire FA_out_1699;
  wire FA_out_1700;
  wire FA_out_1701;
  wire FA_out_1702;
  wire FA_out_1703;
  wire FA_out_1704;
  wire FA_out_1705;
  wire FA_out_1706;
  wire FA_out_1707;
  wire FA_out_1708;
  wire FA_out_1709;
  wire FA_out_1710;
  wire FA_out_1711;
  wire FA_out_1712;
  wire FA_out_1713;
  wire FA_out_1714;
  wire FA_out_1715;
  wire FA_out_1716;
  wire FA_out_1717;
  wire FA_out_1718;
  wire FA_out_1719;
  wire FA_out_1720;
  wire FA_out_1721;
  wire FA_out_1722;
  wire FA_out_1723;
  wire FA_out_1724;
  wire FA_out_1725;
  wire FA_out_1726;
  wire FA_out_1727;
  wire FA_out_1728;
  wire FA_out_1729;
  wire FA_out_1730;
  wire FA_out_1731;
  wire FA_out_1732;
  wire FA_out_1733;
  wire FA_out_1734;
  wire FA_out_1735;
  wire FA_out_1736;
  wire FA_out_1737;
  wire FA_out_1738;
  wire FA_out_1739;
  wire FA_out_1740;
  wire FA_out_1741;
  wire FA_out_1742;
  wire FA_out_1743;
  wire FA_out_1744;
  wire FA_out_1745;
  wire FA_out_1746;
  wire FA_out_1747;
  wire FA_out_1748;
  wire FA_out_1749;
  wire FA_out_1750;
  wire FA_out_1751;
  wire FA_out_1752;
  wire FA_out_1753;
  wire FA_out_1754;
  wire FA_out_1755;
  wire FA_out_1756;
  wire FA_out_1757;
  wire FA_out_1758;
  wire FA_out_1759;
  wire FA_out_1760;
  wire FA_out_1761;
  wire FA_out_1762;
  wire FA_out_1763;
  wire FA_out_1764;
  wire FA_out_1765;
  wire FA_out_1766;
  wire FA_out_1767;
  wire FA_out_1768;
  wire FA_out_1769;
  wire FA_out_1770;
  wire FA_out_1771;
  wire FA_out_1772;
  wire FA_out_1773;
  wire FA_out_1774;
  wire FA_out_1775;
  wire FA_out_1776;
  wire FA_out_1777;
  wire FA_out_1778;
  wire FA_out_1779;
  wire FA_out_1780;
  wire FA_out_1781;
  wire FA_out_1782;
  wire FA_out_1783;
  wire FA_out_1784;
  wire FA_out_1785;
  wire FA_out_1786;
  wire FA_out_1787;
  wire FA_out_1788;
  wire FA_out_1789;
  wire FA_out_1790;
  wire FA_out_1791;
  wire FA_out_1792;
  wire FA_out_1793;
  wire FA_out_1794;
  wire FA_out_1795;
  wire FA_out_1796;
  wire FA_out_1797;
  wire FA_out_1798;
  wire FA_out_1799;
  wire FA_out_1800;
  wire FA_out_1801;
  wire FA_out_1802;
  wire FA_out_1803;
  wire FA_out_1804;
  wire FA_out_1805;
  wire FA_out_1806;
  wire FA_out_1807;
  wire FA_out_1808;
  wire FA_out_1809;
  wire FA_out_1810;
  wire FA_out_1811;
  wire FA_out_1812;
  wire FA_out_1813;
  wire FA_out_1814;
  wire FA_out_1815;
  wire FA_out_1816;
  wire FA_out_1817;
  wire FA_out_1818;
  wire FA_out_1819;
  wire FA_out_1820;
  wire FA_out_1821;
  wire FA_out_1822;
  wire FA_out_1823;
  wire FA_out_1824;
  wire FA_out_1825;
  wire FA_out_1826;
  wire FA_out_1827;
  wire FA_out_1828;
  wire FA_out_1829;
  wire FA_out_1830;
  wire FA_out_1831;
  wire FA_out_1832;
  wire FA_out_1833;
  wire FA_out_1834;
  wire FA_out_1835;
  wire FA_out_1836;
  wire FA_out_1837;
  wire FA_out_1838;
  wire FA_out_1839;
  wire FA_out_1840;
  wire FA_out_1841;
  wire FA_out_1842;
  wire FA_out_1843;
  wire FA_out_1844;
  wire FA_out_1845;
  wire FA_out_1846;
  wire FA_out_1847;
  wire FA_out_1848;
  wire FA_out_1849;
  wire FA_out_1850;
  wire FA_out_1851;
  wire FA_out_1852;
  wire FA_out_1853;
  wire FA_out_1854;
  wire FA_out_1855;
  wire FA_out_1856;
  wire FA_out_1857;
  wire FA_out_1858;
  wire FA_out_1859;
  wire FA_out_1860;
  wire FA_out_1861;
  wire FA_out_1862;
  wire FA_out_1863;
  wire FA_out_1864;
  wire FA_out_1865;
  wire FA_out_1866;
  wire FA_out_1867;
  wire FA_out_1868;
  wire FA_out_1869;
  wire FA_out_1870;
  wire FA_out_1871;
  wire FA_out_1872;
  wire FA_out_1873;
  wire FA_out_1874;
  wire FA_out_1875;
  wire FA_out_1876;
  wire FA_out_1877;
  wire FA_out_1878;
  wire FA_out_1879;
  wire FA_out_1880;
  wire FA_out_1881;
  wire FA_out_1882;
  wire FA_out_1883;
  wire FA_out_1884;
  wire FA_out_1885;
  wire FA_out_1886;
  wire FA_out_1887;
  wire FA_out_1888;
  wire FA_out_1889;
  wire FA_out_1890;
  wire FA_out_1891;
  wire FA_out_1892;
  wire FA_out_1893;
  wire FA_out_1894;
  wire FA_out_1895;
  wire FA_out_1896;
  wire FA_out_1897;
  wire FA_out_1898;
  wire FA_out_1899;
  wire FA_out_1900;
  wire FA_out_1901;
  wire FA_out_1902;
  wire FA_out_1903;
  wire FA_out_1904;
  wire FA_out_1905;
  wire FA_out_1906;
  wire FA_out_1907;
  wire FA_out_1908;
  wire FA_out_1909;
  wire FA_out_1910;
  wire FA_out_1911;
  wire FA_out_1912;
  wire FA_out_1913;
  wire FA_out_1914;
  wire FA_out_1915;
  wire FA_out_1916;
  wire FA_out_1917;
  wire FA_out_1918;
  wire FA_out_1919;
  wire FA_out_1920;
  wire FA_out_1921;
  wire FA_out_1922;
  wire FA_out_1923;
  wire FA_out_1924;
  wire FA_out_1925;
  wire FA_out_1926;
  wire FA_out_1927;
  wire FA_out_1928;
  wire FA_out_1929;
  wire FA_out_1930;
  wire FA_out_1931;
  wire FA_out_1932;
  wire FA_out_1933;
  wire FA_out_1934;
  wire FA_out_1935;
  wire FA_out_1936;
  wire FA_out_1937;
  wire FA_out_1938;
  wire FA_out_1939;
  wire FA_out_1940;
  wire FA_out_1941;
  wire FA_out_1942;
  wire FA_out_1943;
  wire FA_out_1944;
  wire FA_out_1945;
  wire FA_out_1946;
  wire FA_out_1947;
  wire FA_out_1948;
  wire FA_out_1949;
  wire FA_out_1950;
  wire FA_out_1951;
  wire FA_out_1952;
  wire FA_out_1953;
  wire FA_out_1954;
  wire FA_out_1955;
  wire FA_out_1956;
  wire FA_out_1957;
  wire FA_out_1958;
  wire FA_out_1959;
  wire FA_out_1960;
  wire FA_out_1961;
  wire FA_out_1962;
  wire FA_out_1963;
  wire FA_out_1964;
  wire FA_out_1965;
  wire FA_out_1966;
  wire FA_out_1967;
  wire FA_out_1968;
  wire FA_out_1969;
  wire FA_out_1970;
  wire FA_out_1971;
  wire FA_out_1972;
  wire FA_out_1973;
  wire FA_out_1974;
  wire FA_out_1975;
  wire FA_out_1976;
  wire FA_out_1977;
  wire FA_out_1978;
  wire FA_out_1979;
  wire FA_out_1980;
  wire FA_out_1981;
  wire FA_out_1982;
  wire FA_out_1983;
  wire FA_out_1984;
  wire FA_out_1985;
  wire FA_out_1986;
  wire FA_out_1987;
  wire FA_out_1988;
  wire FA_out_1989;
  wire FA_out_1990;
  wire FA_out_1991;
  wire FA_out_1992;
  wire FA_out_1993;
  wire FA_out_1994;
  wire FA_out_1995;
  wire FA_out_1996;
  wire FA_out_1997;
  wire FA_out_1998;
  wire FA_out_1999;
  wire FA_out_2000;
  wire FA_out_2001;
  wire FA_out_2002;
  wire FA_out_2003;
  wire FA_out_2004;
  wire FA_out_2005;
  wire FA_out_2006;
  wire FA_out_2007;
  wire FA_out_2008;
  wire FA_out_2009;
  wire FA_out_2010;
  wire FA_out_2011;
  wire FA_out_2012;
  wire FA_out_2013;
  wire FA_out_2014;
  wire FA_out_2015;
  wire FA_out_2016;
  wire FA_out_2017;
  wire FA_out_2018;
  wire FA_out_2019;
  wire FA_out_2020;
  wire FA_out_2021;
  wire FA_out_2022;
  wire FA_out_2023;
  wire FA_out_2024;
  wire FA_out_2025;
  wire FA_out_2026;
  wire FA_out_2027;
  wire FA_out_2028;
  wire FA_out_2029;
  wire FA_out_2030;
  wire FA_out_2031;
  wire FA_out_2032;
  wire FA_out_2033;
  wire FA_out_2034;
  wire FA_out_2035;
  wire FA_out_2036;
  wire FA_out_2037;
  wire FA_out_2038;
  wire FA_out_2039;
  wire FA_out_2040;
  wire FA_out_2041;
  wire FA_out_2042;
  wire FA_out_2043;
  wire FA_out_2044;
  wire FA_out_2045;
  wire FA_out_2046;
  wire FA_out_2047;
  wire FA_out_2048;
  wire FA_out_2049;
  wire FA_out_2050;
  wire FA_out_2051;
  wire FA_out_2052;
  wire FA_out_2053;
  wire FA_out_2054;
  wire FA_out_2055;
  wire FA_out_2056;
  wire FA_out_2057;
  wire FA_out_2058;
  wire FA_out_2059;
  wire FA_out_2060;
  wire FA_out_2061;
  wire FA_out_2062;
  wire FA_out_2063;
  wire FA_out_2064;
  wire FA_out_2065;
  wire FA_out_2066;
  wire FA_out_2067;
  wire FA_out_2068;
  wire FA_out_2069;
  wire FA_out_2070;
  wire FA_out_2071;
  wire FA_out_2072;
  wire FA_out_2073;
  wire FA_out_2074;
  wire FA_out_2075;
  wire FA_out_2076;
  wire FA_out_2077;
  wire FA_out_2078;
  wire FA_out_2079;
  wire FA_out_2080;
  wire FA_out_2081;
  wire FA_out_2082;
  wire FA_out_2083;
  wire FA_out_2084;
  wire FA_out_2085;
  wire FA_out_2086;
  wire FA_out_2087;
  wire FA_out_2088;
  wire FA_out_2089;
  wire FA_out_2090;
  wire FA_out_2091;
  wire FA_out_2092;
  wire FA_out_2093;
  wire FA_out_2094;
  wire FA_out_2095;
  wire FA_out_2096;
  wire FA_out_2097;
  wire FA_out_2098;
  wire FA_out_2099;
  wire FA_out_2100;
  wire FA_out_2101;
  wire FA_out_2102;
  wire FA_out_2103;
  wire FA_out_2104;
  wire FA_out_2105;
  wire FA_out_2106;
  wire FA_out_2107;
  wire FA_out_2108;
  wire FA_out_2109;
  wire FA_out_2110;
  wire FA_out_2111;
  wire FA_out_2112;
  wire FA_out_2113;
  wire FA_out_2114;
  wire FA_out_2115;
  wire FA_out_2116;
  wire FA_out_2117;
  wire FA_out_2118;
  wire FA_out_2119;
  wire FA_out_2120;
  wire FA_out_2121;
  wire FA_out_2122;
  wire FA_out_2123;
  wire FA_out_2124;
  wire FA_out_2125;
  wire FA_out_2126;
  wire FA_out_2127;
  wire FA_out_2128;
  wire FA_out_2129;
  wire FA_out_2130;
  wire FA_out_2131;
  wire FA_out_2132;
  wire FA_out_2133;
  wire FA_out_2134;
  wire FA_out_2135;
  wire FA_out_2136;
  wire FA_out_2137;
  wire FA_out_2138;
  wire FA_out_2139;
  wire FA_out_2140;
  wire FA_out_2141;
  wire FA_out_2142;
  wire FA_out_2143;
  wire FA_out_2144;
  wire FA_out_2145;
  wire FA_out_2146;
  wire FA_out_2147;
  wire FA_out_2148;
  wire FA_out_2149;
  wire FA_out_2150;
  wire FA_out_2151;
  wire FA_out_2152;
  wire FA_out_2153;
  wire FA_out_2154;
  wire FA_out_2155;
  wire FA_out_2156;
  wire FA_out_2157;
  wire FA_out_2158;
  wire FA_out_2159;
  wire FA_out_2160;
  wire FA_out_2161;
  wire FA_out_2162;
  wire FA_out_2163;
  wire FA_out_2164;
  wire FA_out_2165;
  wire FA_out_2166;
  wire FA_out_2167;
  wire FA_out_2168;
  wire FA_out_2169;
  wire FA_out_2170;
  wire FA_out_2171;
  wire FA_out_2172;
  wire FA_out_2173;
  wire FA_out_2174;
  wire FA_out_2175;
  wire FA_out_2176;
  wire FA_out_2177;
  wire FA_out_2178;
  wire FA_out_2179;
  wire FA_out_2180;
  wire FA_out_2181;
  wire FA_out_2182;
  wire FA_out_2183;
  wire FA_out_2184;
  wire FA_out_2185;
  wire FA_out_2186;
  wire FA_out_2187;
  wire FA_out_2188;
  wire FA_out_2189;
  wire FA_out_2190;
  wire FA_out_2191;
  wire FA_out_2192;
  wire FA_out_2193;
  wire FA_out_2194;
  wire FA_out_2195;
  wire FA_out_2196;
  wire FA_out_2197;
  wire FA_out_2198;
  wire FA_out_2199;
  wire FA_out_2200;
  wire FA_out_2201;
  wire FA_out_2202;
  wire FA_out_2203;
  wire FA_out_2204;
  wire FA_out_2205;
  wire FA_out_2206;
  wire FA_out_2207;
  wire FA_out_2208;
  wire FA_out_2209;
  wire FA_out_2210;
  wire FA_out_2211;
  wire FA_out_2212;
  wire FA_out_2213;
  wire FA_out_2214;
  wire FA_out_2215;
  wire FA_out_2216;
  wire FA_out_2217;
  wire FA_out_2218;
  wire FA_out_2219;
  wire FA_out_2220;
  wire FA_out_2221;
  wire FA_out_2222;
  wire FA_out_2223;
  wire FA_out_2224;
  wire FA_out_2225;
  wire FA_out_2226;
  wire FA_out_2227;
  wire FA_out_2228;
  wire FA_out_2229;
  wire FA_out_2230;
  wire FA_out_2231;
  wire FA_out_2232;
  wire FA_out_2233;
  wire FA_out_2234;
  wire FA_out_2235;
  wire FA_out_2236;
  wire FA_out_2237;
  wire FA_out_2238;
  wire FA_out_2239;
  wire FA_out_2240;
  wire FA_out_2241;
  wire FA_out_2242;
  wire FA_out_2243;
  wire FA_out_2244;
  wire FA_out_2245;
  wire FA_out_2246;
  wire FA_out_2247;
  wire FA_out_2248;
  wire FA_out_2249;
  wire FA_out_2250;
  wire FA_out_2251;
  wire FA_out_2252;
  wire FA_out_2253;
  wire FA_out_2254;
  wire FA_out_2255;
  wire FA_out_2256;
  wire FA_out_2257;
  wire FA_out_2258;
  wire FA_out_2259;
  wire FA_out_2260;
  wire FA_out_2261;
  wire FA_out_2262;
  wire FA_out_2263;
  wire FA_out_2264;
  wire FA_out_2265;
  wire FA_out_2266;
  wire FA_out_2267;
  wire FA_out_2268;
  wire FA_out_2269;
  wire FA_out_2270;
  wire FA_out_2271;
  wire FA_out_2272;
  wire FA_out_2273;
  wire FA_out_2274;
  wire FA_out_2275;
  wire FA_out_2276;
  wire FA_out_2277;
  wire FA_out_2278;
  wire FA_out_2279;
  wire FA_out_2280;
  wire FA_out_2281;
  wire FA_out_2282;
  wire FA_out_2283;
  wire FA_out_2284;
  wire FA_out_2285;
  wire FA_out_2286;
  wire FA_out_2287;
  wire FA_out_2288;
  wire FA_out_2289;
  wire FA_out_2290;
  wire FA_out_2291;
  wire FA_out_2292;
  wire FA_out_2293;
  wire FA_out_2294;
  wire FA_out_2295;
  wire FA_out_2296;
  wire FA_out_2297;
  wire FA_out_2298;
  wire FA_out_2299;
  wire FA_out_2300;
  wire FA_out_2301;
  wire FA_out_2302;
  wire FA_out_2303;
  wire FA_out_2304;
  wire FA_out_2305;
  wire FA_out_2306;
  wire FA_out_2307;
  wire FA_out_2308;
  wire FA_out_2309;
  wire FA_out_2310;
  wire FA_out_2311;
  wire FA_out_2312;
  wire FA_out_2313;
  wire FA_out_2314;
  wire FA_out_2315;
  wire FA_out_2316;
  wire FA_out_2317;
  wire FA_out_2318;
  wire FA_out_2319;
  wire FA_out_2320;
  wire FA_out_2321;
  wire FA_out_2322;
  wire FA_out_2323;
  wire FA_out_2324;
  wire FA_out_2325;
  wire FA_out_2326;
  wire FA_out_2327;
  wire FA_out_2328;
  wire FA_out_2329;
  wire FA_out_2330;
  wire FA_out_2331;
  wire FA_out_2332;
  wire FA_out_2333;
  wire FA_out_2334;
  wire FA_out_2335;
  wire FA_out_2336;
  wire FA_out_2337;
  wire FA_out_2338;
  wire FA_out_2339;
  wire FA_out_2340;
  wire FA_out_2341;
  wire FA_out_2342;
  wire FA_out_2343;
  wire FA_out_2344;
  wire FA_out_2345;
  wire FA_out_2346;
  wire FA_out_2347;
  wire FA_out_2348;
  wire FA_out_2349;
  wire FA_out_2350;
  wire FA_out_2351;
  wire FA_out_2352;
  wire FA_out_2353;
  wire FA_out_2354;
  wire FA_out_2355;
  wire FA_out_2356;
  wire FA_out_2357;
  wire FA_out_2358;
  wire FA_out_2359;
  wire FA_out_2360;
  wire FA_out_2361;
  wire FA_out_2362;
  wire FA_out_2363;
  wire FA_out_2364;
  wire FA_out_2365;
  wire FA_out_2366;
  wire FA_out_2367;
  wire FA_out_2368;
  wire FA_out_2369;
  wire FA_out_2370;
  wire FA_out_2371;
  wire FA_out_2372;
  wire FA_out_2373;
  wire FA_out_2374;
  wire FA_out_2375;
  wire FA_out_2376;
  wire FA_out_2377;
  wire FA_out_2378;
  wire FA_out_2379;
  wire FA_out_2380;
  wire FA_out_2381;
  wire FA_out_2382;
  wire FA_out_2383;
  wire FA_out_2384;
  wire FA_out_2385;
  wire FA_out_2386;
  wire FA_out_2387;
  wire FA_out_2388;
  wire FA_out_2389;
  wire FA_out_2390;
  wire FA_out_2391;
  wire FA_out_2392;
  wire FA_out_2393;
  wire FA_out_2394;
  wire FA_out_2395;
  wire FA_out_2396;
  wire FA_out_2397;
  wire FA_out_2398;
  wire FA_out_2399;
  wire FA_out_2400;
  wire FA_out_2401;
  wire FA_out_2402;
  wire FA_out_2403;
  wire FA_out_2404;
  wire FA_out_2405;
  wire FA_out_2406;
  wire FA_out_2407;
  wire FA_out_2408;
  wire FA_out_2409;
  wire FA_out_2410;
  wire FA_out_2411;
  wire FA_out_2412;
  wire FA_out_2413;
  wire FA_out_2414;
  wire FA_out_2415;
  wire FA_out_2416;
  wire FA_out_2417;
  wire FA_out_2418;
  wire FA_out_2419;
  wire FA_out_2420;
  wire FA_out_2421;
  wire FA_out_2422;
  wire FA_out_2423;
  wire FA_out_2424;
  wire FA_out_2425;
  wire FA_out_2426;
  wire FA_out_2427;
  wire FA_out_2428;
  wire FA_out_2429;
  wire FA_out_2430;
  wire FA_out_2431;
  wire FA_out_2432;
  wire FA_out_2433;
  wire FA_out_2434;
  wire FA_out_2435;
  wire FA_out_2436;
  wire FA_out_2437;
  wire FA_out_2438;
  wire FA_out_2439;
  wire FA_out_2440;
  wire FA_out_2441;
  wire FA_out_2442;
  wire FA_out_2443;
  wire FA_out_2444;
  wire FA_out_2445;
  wire FA_out_2446;
  wire FA_out_2447;
  wire FA_out_2448;
  wire FA_out_2449;
  wire FA_out_2450;
  wire FA_out_2451;
  wire FA_out_2452;
  wire FA_out_2453;
  wire FA_out_2454;
  wire FA_out_2455;
  wire FA_out_2456;
  wire FA_out_2457;
  wire FA_out_2458;
  wire FA_out_2459;
  wire FA_out_2460;
  wire FA_out_2461;
  wire FA_out_2462;
  wire FA_out_2463;
  wire FA_out_2464;
  wire FA_out_2465;
  wire FA_out_2466;
  wire FA_out_2467;
  wire FA_out_2468;
  wire FA_out_2469;
  wire FA_out_2470;
  wire FA_out_2471;
  wire FA_out_2472;
  wire FA_out_2473;
  wire FA_out_2474;
  wire FA_out_2475;
  wire FA_out_2476;
  wire FA_out_2477;
  wire FA_out_2478;
  wire FA_out_2479;
  wire FA_out_2480;
  wire FA_out_2481;
  wire FA_out_2482;
  wire FA_out_2483;
  wire FA_out_2484;
  wire FA_out_2485;
  wire FA_out_2486;
  wire FA_out_2487;
  wire FA_out_2488;
  wire FA_out_2489;
  wire FA_out_2490;
  wire FA_out_2491;
  wire FA_out_2492;
  wire FA_out_2493;
  wire FA_out_2494;
  wire FA_out_2495;
  wire FA_out_2496;
  wire FA_out_2497;
  wire FA_out_2498;
  wire FA_out_2499;
  wire FA_out_2500;
  wire FA_out_2501;
  wire FA_out_2502;
  wire FA_out_2503;
  wire FA_out_2504;
  wire FA_out_2505;
  wire FA_out_2506;
  wire FA_out_2507;
  wire FA_out_2508;
  wire FA_out_2509;
  wire FA_out_2510;
  wire FA_out_2511;
  wire FA_out_2512;
  wire FA_out_2513;
  wire FA_out_2514;
  wire FA_out_2515;
  wire FA_out_2516;
  wire FA_out_2517;
  wire FA_out_2518;
  wire FA_out_2519;
  wire FA_out_2520;
  wire FA_out_2521;
  wire FA_out_2522;
  wire FA_out_2523;
  wire FA_out_2524;
  wire FA_out_2525;
  wire FA_out_2526;
  wire FA_out_2527;
  wire FA_out_2528;
  wire FA_out_2529;
  wire FA_out_2530;
  wire FA_out_2531;
  wire FA_out_2532;
  wire FA_out_2533;
  wire FA_out_2534;
  wire FA_out_2535;
  wire FA_out_2536;
  wire FA_out_2537;
  wire FA_out_2538;
  wire FA_out_2539;
  wire FA_out_2540;
  wire FA_out_2541;
  wire FA_out_2542;
  wire FA_out_2543;
  wire FA_out_2544;
  wire FA_out_2545;
  wire FA_out_2546;
  wire FA_out_2547;
  wire FA_out_2548;
  wire FA_out_2549;
  wire FA_out_2550;
  wire FA_out_2551;
  wire FA_out_2552;
  wire FA_out_2553;
  wire FA_out_2554;
  wire FA_out_2555;
  wire FA_out_2556;
  wire FA_out_2557;
  wire FA_out_2558;
  wire FA_out_2559;
  wire FA_out_2560;
  wire FA_out_2561;
  wire FA_out_2562;
  wire FA_out_2563;
  wire FA_out_2564;
  wire FA_out_2565;
  wire FA_out_2566;
  wire FA_out_2567;
  wire FA_out_2568;
  wire FA_out_2569;
  wire FA_out_2570;
  wire FA_out_2571;
  wire FA_out_2572;
  wire FA_out_2573;
  wire FA_out_2574;
  wire FA_out_2575;
  wire FA_out_2576;
  wire FA_out_2577;
  wire FA_out_2578;
  wire FA_out_2579;
  wire FA_out_2580;
  wire FA_out_2581;
  wire FA_out_2582;
  wire FA_out_2583;
  wire FA_out_2584;
  wire FA_out_2585;
  wire FA_out_2586;
  wire FA_out_2587;
  wire FA_out_2588;
  wire FA_out_2589;
  wire FA_out_2590;
  wire FA_out_2591;
  wire FA_out_2592;
  wire FA_out_2593;
  wire FA_out_2594;
  wire FA_out_2595;
  wire FA_out_2596;
  wire FA_out_2597;
  wire FA_out_2598;
  wire FA_out_2599;
  wire FA_out_2600;
  wire FA_out_2601;
  wire FA_out_2602;
  wire FA_out_2603;
  wire FA_out_2604;
  wire FA_out_2605;
  wire FA_out_2606;
  wire FA_out_2607;
  wire FA_out_2608;
  wire FA_out_2609;
  wire FA_out_2610;
  wire FA_out_2611;
  wire FA_out_2612;
  wire FA_out_2613;
  wire FA_out_2614;
  wire FA_out_2615;
  wire FA_out_2616;
  wire FA_out_2617;
  wire FA_out_2618;
  wire FA_out_2619;
  wire FA_out_2620;
  wire FA_out_2621;
  wire FA_out_2622;
  wire FA_out_2623;
  wire FA_out_2624;
  wire FA_out_2625;
  wire FA_out_2626;
  wire FA_out_2627;
  wire FA_out_2628;
  wire FA_out_2629;
  wire FA_out_2630;
  wire FA_out_2631;
  wire FA_out_2632;
  wire FA_out_2633;
  wire FA_out_2634;
  wire FA_out_2635;
  wire FA_out_2636;
  wire FA_out_2637;
  wire FA_out_2638;
  wire FA_out_2639;
  wire FA_out_2640;
  wire FA_out_2641;
  wire FA_out_2642;
  wire FA_out_2643;
  wire FA_out_2644;
  wire FA_out_2645;
  wire FA_out_2646;
  wire FA_out_2647;
  wire FA_out_2648;
  wire FA_out_2649;
  wire FA_out_2650;
  wire FA_out_2651;
  wire FA_out_2652;
  wire FA_out_2653;
  wire FA_out_2654;
  wire FA_out_2655;
  wire FA_out_2656;
  wire FA_out_2657;
  wire FA_out_2658;
  wire FA_out_2659;
  wire FA_out_2660;
  wire FA_out_2661;
  wire FA_out_2662;
  wire FA_out_2663;
  wire FA_out_2664;
  wire FA_out_2665;
  wire FA_out_2666;
  wire FA_out_2667;
  wire FA_out_2668;
  wire FA_out_2669;
  wire FA_out_2670;
  wire FA_out_2671;
  wire FA_out_2672;
  wire FA_out_2673;
  wire FA_out_2674;
  wire FA_out_2675;
  wire FA_out_2676;
  wire FA_out_2677;
  wire FA_out_2678;
  wire FA_out_2679;
  wire FA_out_2680;
  wire FA_out_2681;
  wire FA_out_2682;
  wire FA_out_2683;
  wire FA_out_2684;
  wire FA_out_2685;
  wire FA_out_2686;
  wire FA_out_2687;
  wire FA_out_2688;
  wire FA_out_2689;
  wire FA_out_2690;
  wire FA_out_2691;
  wire FA_out_2692;
  wire FA_out_2693;
  wire FA_out_2694;
  wire FA_out_2695;
  wire FA_out_2696;
  wire FA_out_2697;
  wire FA_out_2698;
  wire FA_out_2699;
  wire FA_out_2700;
  wire FA_out_2701;
  wire FA_out_2702;
  wire FA_out_2703;
  wire FA_out_2704;
  wire FA_out_2705;
  wire FA_out_2706;
  wire FA_out_2707;
  wire FA_out_2708;
  wire FA_out_2709;
  wire FA_out_2710;
  wire FA_out_2711;
  wire FA_out_2712;
  wire FA_out_2713;
  wire FA_out_2714;
  wire FA_out_2715;
  wire FA_out_2716;
  wire FA_out_2717;
  wire FA_out_2718;
  wire FA_out_2719;
  wire FA_out_2720;
  wire FA_out_2721;
  wire FA_out_2722;
  wire FA_out_2723;
  wire FA_out_2724;
  wire FA_out_2725;
  wire FA_out_2726;
  wire FA_out_2727;
  wire FA_out_2728;
  wire FA_out_2729;
  wire FA_out_2730;
  wire FA_out_2731;
  wire FA_out_2732;
  wire FA_out_2733;
  wire FA_out_2734;
  wire FA_out_2735;
  wire FA_out_2736;
  wire FA_out_2737;
  wire FA_out_2738;
  wire FA_out_2739;
  wire FA_out_2740;
  wire FA_out_2741;
  wire FA_out_2742;
  wire FA_out_2743;
  wire FA_out_2744;
  wire FA_out_2745;
  wire FA_out_2746;
  wire FA_out_2747;
  wire FA_out_2748;
  wire FA_out_2749;
  wire FA_out_2750;
  wire FA_out_2751;
  wire FA_out_2752;
  wire FA_out_2753;
  wire FA_out_2754;
  wire FA_out_2755;
  wire FA_out_2756;
  wire FA_out_2757;
  wire FA_out_2758;
  wire FA_out_2759;
  wire FA_out_2760;
  wire FA_out_2761;
  wire FA_out_2762;
  wire FA_out_2763;
  wire FA_out_2764;
  wire FA_out_2765;
  wire FA_out_2766;
  wire FA_out_2767;
  wire FA_out_2768;
  wire FA_out_2769;
  wire FA_out_2770;
  wire FA_out_2771;
  wire FA_out_2772;
  wire FA_out_2773;
  wire FA_out_2774;
  wire FA_out_2775;
  wire FA_out_2776;
  wire FA_out_2777;
  wire FA_out_2778;
  wire FA_out_2779;
  wire FA_out_2780;
  wire FA_out_2781;
  wire FA_out_2782;
  wire FA_out_2783;
  wire FA_out_2784;
  wire FA_out_2785;
  wire FA_out_2786;
  wire FA_out_2787;
  wire FA_out_2788;
  wire FA_out_2789;
  wire FA_out_2790;
  wire FA_out_2791;
  wire FA_out_2792;
  wire FA_out_2793;
  wire FA_out_2794;
  wire FA_out_2795;
  wire FA_out_2796;
  wire FA_out_2797;
  wire FA_out_2798;
  wire FA_out_2799;
  wire FA_out_2800;
  wire FA_out_2801;
  wire FA_out_2802;
  wire FA_out_2803;
  wire FA_out_2804;
  wire FA_out_2805;
  wire FA_out_2806;
  wire FA_out_2807;
  wire FA_out_2808;
  wire FA_out_2809;
  wire FA_out_2810;
  wire FA_out_2811;
  wire FA_out_2812;
  wire FA_out_2813;
  wire FA_out_2814;
  wire FA_out_2815;
  wire FA_out_2816;
  wire FA_out_2817;
  wire FA_out_2818;
  wire FA_out_2819;
  wire FA_out_2820;
  wire FA_out_2821;
  wire FA_out_2822;
  wire FA_out_2823;
  wire FA_out_2824;
  wire FA_out_2825;
  wire FA_out_2826;
  wire FA_out_2827;
  wire FA_out_2828;
  wire FA_out_2829;
  wire FA_out_2830;
  wire FA_out_2831;
  wire FA_out_2832;
  wire FA_out_2833;
  wire FA_out_2834;
  wire FA_out_2835;
  wire FA_out_2836;
  wire FA_out_2837;
  wire FA_out_2838;
  wire FA_out_2839;
  wire FA_out_2840;
  wire FA_out_2841;
  wire FA_out_2842;
  wire FA_out_2843;
  wire FA_out_2844;
  wire FA_out_2845;
  wire FA_out_2846;
  wire FA_out_2847;
  wire FA_out_2848;
  wire FA_out_2849;
  wire FA_out_2850;
  wire FA_out_2851;
  wire FA_out_2852;
  wire FA_out_2853;
  wire FA_out_2854;
  wire FA_out_2855;
  wire FA_out_2856;
  wire FA_out_2857;
  wire FA_out_2858;
  wire FA_out_2859;
  wire FA_out_2860;
  wire FA_out_2861;
  wire FA_out_2862;
  wire FA_out_2863;
  wire FA_out_2864;
  wire FA_out_2865;
  wire FA_out_2866;
  wire FA_out_2867;
  wire FA_out_2868;
  wire FA_out_2869;
  wire FA_out_2870;
  wire FA_out_2871;
  wire FA_out_2872;
  wire FA_out_2873;
  wire FA_out_2874;
  wire FA_out_2875;
  wire FA_out_2876;
  wire FA_out_2877;
  wire FA_out_2878;
  wire FA_out_2879;
  wire FA_out_2880;
  wire FA_out_2881;
  wire FA_out_2882;
  wire FA_out_2883;
  wire FA_out_2884;
  wire FA_out_2885;
  wire FA_out_2886;
  wire FA_out_2887;
  wire FA_out_2888;
  wire FA_out_2889;
  wire FA_out_2890;
  wire FA_out_2891;
  wire FA_out_2892;
  wire FA_out_2893;
  wire FA_out_2894;
  wire FA_out_2895;
  wire FA_out_2896;
  wire FA_out_2897;
  wire FA_out_2898;
  wire FA_out_2899;
  wire FA_out_2900;
  wire FA_out_2901;
  wire FA_out_2902;
  wire FA_out_2903;
  wire FA_out_2904;
  wire FA_out_2905;
  wire FA_out_2906;
  wire FA_out_2907;
  wire FA_out_2908;
  wire FA_out_2909;
  wire FA_out_2910;
  wire FA_out_2911;
  wire FA_out_2912;
  wire FA_out_2913;
  wire FA_out_2914;
  wire FA_out_2915;
  wire FA_out_2916;
  wire FA_out_2917;
  wire FA_out_2918;
  wire FA_out_2919;
  wire FA_out_2920;
  wire FA_out_2921;
  wire FA_out_2922;
  wire FA_out_2923;
  wire FA_out_2924;
  wire FA_out_2925;
  wire FA_out_2926;
  wire FA_out_2927;
  wire FA_out_2928;
  wire FA_out_2929;
  wire FA_out_2930;
  wire FA_out_2931;
  wire FA_out_2932;
  wire FA_out_2933;
  wire FA_out_2934;
  wire FA_out_2935;
  wire FA_out_2936;
  wire FA_out_2937;
  wire FA_out_2938;
  wire FA_out_2939;
  wire FA_out_2940;
  wire FA_out_2941;
  wire FA_out_2942;
  wire FA_out_2943;
  wire FA_out_2944;
  wire FA_out_2945;
  wire FA_out_2946;
  wire FA_out_2947;
  wire FA_out_2948;
  wire FA_out_2949;
  wire FA_out_2950;
  wire FA_out_2951;
  wire FA_out_2952;
  wire FA_out_2953;
  wire FA_out_2954;
  wire FA_out_2955;
  wire FA_out_2956;
  wire FA_out_2957;
  wire FA_out_2958;
  wire FA_out_2959;
  wire FA_out_2960;
  wire FA_out_2961;
  wire FA_out_2962;
  wire FA_out_2963;
  wire FA_out_2964;
  wire FA_out_2965;
  wire FA_out_2966;
  wire FA_out_2967;
  wire FA_out_2968;
  wire FA_out_2969;
  wire FA_out_2970;
  wire FA_out_2971;
  wire FA_out_2972;
  wire FA_out_2973;
  wire FA_out_2974;
  wire FA_out_2975;
  wire FA_out_2976;
  wire FA_out_2977;
  wire FA_out_2978;
  wire FA_out_2979;
  wire FA_out_2980;
  wire FA_out_2981;
  wire FA_out_2982;
  wire FA_out_2983;
  wire FA_out_2984;
  wire FA_out_2985;
  wire FA_out_2986;
  wire FA_out_2987;
  wire FA_out_2988;
  wire FA_out_2989;
  wire FA_out_2990;
  wire FA_out_2991;
  wire FA_out_2992;
  wire FA_out_2993;
  wire FA_out_2994;
  wire FA_out_2995;
  wire FA_out_2996;
  wire FA_out_2997;
  wire FA_out_2998;
  wire FA_out_2999;
  wire FA_out_3000;
  wire FA_out_3001;
  wire FA_out_3002;
  wire FA_out_3003;
  wire FA_out_3004;
  wire FA_out_3005;
  wire FA_out_3006;
  wire FA_out_3007;
  wire FA_out_3008;
  wire FA_out_3009;
  wire FA_out_3010;
  wire FA_out_3011;
  wire FA_out_3012;
  wire FA_out_3013;
  wire FA_out_3014;
  wire FA_out_3015;
  wire FA_out_3016;
  wire FA_out_3017;
  wire FA_out_3018;
  wire FA_out_3019;
  wire FA_out_3020;
  wire FA_out_3021;
  wire FA_out_3022;
  wire FA_out_3023;
  wire FA_out_3024;
  wire FA_out_3025;
  wire FA_out_3026;
  wire FA_out_3027;
  wire FA_out_3028;
  wire FA_out_3029;
  wire FA_out_3030;
  wire FA_out_3031;
  wire FA_out_3032;
  wire FA_out_3033;
  wire FA_out_3034;
  wire FA_out_3035;
  wire FA_out_3036;
  wire FA_out_3037;
  wire FA_out_3038;
  wire FA_out_3039;
  wire FA_out_3040;
  wire FA_out_3041;
  wire FA_out_3042;
  wire FA_out_3043;
  wire FA_out_3044;
  wire FA_out_3045;
  wire FA_out_3046;
  wire FA_out_3047;
  wire FA_out_3048;
  wire FA_out_3049;
  wire FA_out_3050;
  wire FA_out_3051;
  wire FA_out_3052;
  wire FA_out_3053;
  wire FA_out_3054;
  wire FA_out_3055;
  wire FA_out_3056;
  wire FA_out_3057;
  wire FA_out_3058;
  wire FA_out_3059;
  wire FA_out_3060;
  wire FA_out_3061;
  wire FA_out_3062;
  wire FA_out_3063;
  wire FA_out_3064;
  wire FA_out_3065;
  wire FA_out_3066;
  wire FA_out_3067;
  wire FA_out_3068;
  wire FA_out_3069;
  wire FA_out_3070;
  wire FA_out_3071;
  wire FA_out_3072;
  wire FA_out_3073;
  wire FA_out_3074;
  wire FA_out_3075;
  wire FA_out_3076;
  wire FA_out_3077;
  wire FA_out_3078;
  wire FA_out_3079;
  wire FA_out_3080;
  wire FA_out_3081;
  wire FA_out_3082;
  wire FA_out_3083;
  wire FA_out_3084;
  wire FA_out_3085;
  wire FA_out_3086;
  wire FA_out_3087;
  wire FA_out_3088;
  wire FA_out_3089;
  wire FA_out_3090;
  wire FA_out_3091;
  wire FA_out_3092;
  wire FA_out_3093;
  wire FA_out_3094;
  wire FA_out_3095;
  wire FA_out_3096;
  wire FA_out_3097;
  wire FA_out_3098;
  wire FA_out_3099;
  wire FA_out_3100;
  wire FA_out_3101;
  wire FA_out_3102;
  wire FA_out_3103;
  wire FA_out_3104;
  wire FA_out_3105;
  wire FA_out_3106;
  wire FA_out_3107;
  wire FA_out_3108;
  wire FA_out_3109;
  wire FA_out_3110;
  wire FA_out_3111;
  wire FA_out_3112;
  wire FA_out_3113;
  wire FA_out_3114;
  wire FA_out_3115;
  wire FA_out_3116;
  wire FA_out_3117;
  wire FA_out_3118;
  wire FA_out_3119;
  wire FA_out_3120;
  wire FA_out_3121;
  wire FA_out_3122;
  wire FA_out_3123;
  wire FA_out_3124;
  wire FA_out_3125;
  wire FA_out_3126;
  wire FA_out_3127;
  wire FA_out_3128;
  wire FA_out_3129;
  wire FA_out_3130;
  wire FA_out_3131;
  wire FA_out_3132;
  wire FA_out_3133;
  wire FA_out_3134;
  wire FA_out_3135;
  wire FA_out_3136;
  wire FA_out_3137;
  wire FA_out_3138;
  wire FA_out_3139;
  wire FA_out_3140;
  wire FA_out_3141;
  wire FA_out_3142;
  wire FA_out_3143;
  wire FA_out_3144;
  wire FA_out_3145;
  wire FA_out_3146;
  wire FA_out_3147;
  wire FA_out_3148;
  wire FA_out_3149;
  wire FA_out_3150;
  wire FA_out_3151;
  wire FA_out_3152;
  wire FA_out_3153;
  wire FA_out_3154;
  wire FA_out_3155;
  wire FA_out_3156;
  wire FA_out_3157;
  wire FA_out_3158;
  wire FA_out_3159;
  wire FA_out_3160;
  wire FA_out_3161;
  wire FA_out_3162;
  wire FA_out_3163;
  wire FA_out_3164;
  wire FA_out_3165;
  wire FA_out_3166;
  wire FA_out_3167;
  wire FA_out_3168;
  wire FA_out_3169;
  wire FA_out_3170;
  wire FA_out_3171;
  wire FA_out_3172;
  wire FA_out_3173;
  wire FA_out_3174;
  wire FA_out_3175;
  wire FA_out_3176;
  wire FA_out_3177;
  wire FA_out_3178;
  wire FA_out_3179;
  wire FA_out_3180;
  wire FA_out_3181;
  wire FA_out_3182;
  wire FA_out_3183;
  wire FA_out_3184;
  wire FA_out_3185;
  wire FA_out_3186;
  wire FA_out_3187;
  wire FA_out_3188;
  wire FA_out_3189;
  wire FA_out_3190;
  wire FA_out_3191;
  wire FA_out_3192;
  wire FA_out_3193;
  wire FA_out_3194;
  wire FA_out_3195;
  wire FA_out_3196;
  wire FA_out_3197;
  wire FA_out_3198;
  wire FA_out_3199;
  wire FA_out_3200;
  wire FA_out_3201;
  wire FA_out_3202;
  wire FA_out_3203;
  wire FA_out_3204;
  wire FA_out_3205;
  wire FA_out_3206;
  wire FA_out_3207;
  wire FA_out_3208;
  wire FA_out_3209;
  wire FA_out_3210;
  wire FA_out_3211;
  wire FA_out_3212;
  wire FA_out_3213;
  wire FA_out_3214;
  wire FA_out_3215;
  wire FA_out_3216;
  wire FA_out_3217;
  wire FA_out_3218;
  wire FA_out_3219;
  wire FA_out_3220;
  wire FA_out_3221;
  wire FA_out_3222;
  wire FA_out_3223;
  wire FA_out_3224;
  wire FA_out_3225;
  wire FA_out_3226;
  wire FA_out_3227;
  wire FA_out_3228;
  wire FA_out_3229;
  wire FA_out_3230;
  wire FA_out_3231;
  wire FA_out_3232;
  wire FA_out_3233;
  wire FA_out_3234;
  wire FA_out_3235;
  wire FA_out_3236;
  wire FA_out_3237;
  wire FA_out_3238;
  wire FA_out_3239;
  wire FA_out_3240;
  wire FA_out_3241;
  wire FA_out_3242;
  wire FA_out_3243;
  wire FA_out_3244;
  wire FA_out_3245;
  wire FA_out_3246;
  wire FA_out_3247;
  wire FA_out_3248;
  wire FA_out_3249;
  wire FA_out_3250;
  wire FA_out_3251;
  wire FA_out_3252;
  wire FA_out_3253;
  wire FA_out_3254;
  wire FA_out_3255;
  wire FA_out_3256;
  wire FA_out_3257;
  wire FA_out_3258;
  wire FA_out_3259;
  wire FA_out_3260;
  wire FA_out_3261;
  wire FA_out_3262;
  wire FA_out_3263;
  wire FA_out_3264;
  wire FA_out_3265;
  wire FA_out_3266;
  wire FA_out_3267;
  wire FA_out_3268;
  wire FA_out_3269;
  wire FA_out_3270;
  wire FA_out_3271;
  wire FA_out_3272;
  wire FA_out_3273;
  wire FA_out_3274;
  wire FA_out_3275;
  wire FA_out_3276;
  wire FA_out_3277;
  wire FA_out_3278;
  wire FA_out_3279;
  wire FA_out_3280;
  wire FA_out_3281;
  wire FA_out_3282;
  wire FA_out_3283;
  wire FA_out_3284;
  wire FA_out_3285;
  wire FA_out_3286;
  wire FA_out_3287;
  wire FA_out_3288;
  wire FA_out_3289;
  wire FA_out_3290;
  wire FA_out_3291;
  wire FA_out_3292;
  wire FA_out_3293;
  wire FA_out_3294;
  wire FA_out_3295;
  wire FA_out_3296;
  wire FA_out_3297;
  wire FA_out_3298;
  wire FA_out_3299;
  wire FA_out_3300;
  wire FA_out_3301;
  wire FA_out_3302;
  wire FA_out_3303;
  wire FA_out_3304;
  wire FA_out_3305;
  wire FA_out_3306;
  wire FA_out_3307;
  wire FA_out_3308;
  wire FA_out_3309;
  wire FA_out_3310;
  wire FA_out_3311;
  wire FA_out_3312;
  wire FA_out_3313;
  wire FA_out_3314;
  wire FA_out_3315;
  wire FA_out_3316;
  wire FA_out_3317;
  wire FA_out_3318;
  wire FA_out_3319;
  wire FA_out_3320;
  wire FA_out_3321;
  wire FA_out_3322;
  wire FA_out_3323;
  wire FA_out_3324;
  wire FA_out_3325;
  wire FA_out_3326;
  wire FA_out_3327;
  wire FA_out_3328;
  wire FA_out_3329;
  wire FA_out_3330;
  wire FA_out_3331;
  wire FA_out_3332;
  wire FA_out_3333;
  wire FA_out_3334;
  wire FA_out_3335;
  wire FA_out_3336;
  wire FA_out_3337;
  wire FA_out_3338;
  wire FA_out_3339;
  wire FA_out_3340;
  wire FA_out_3341;
  wire FA_out_3342;
  wire FA_out_3343;
  wire FA_out_3344;
  wire FA_out_3345;
  wire FA_out_3346;
  wire FA_out_3347;
  wire FA_out_3348;
  wire FA_out_3349;
  wire FA_out_3350;
  wire FA_out_3351;
  wire FA_out_3352;
  wire FA_out_3353;
  wire FA_out_3354;
  wire FA_out_3355;
  wire FA_out_3356;
  wire FA_out_3357;
  wire FA_out_3358;
  wire FA_out_3359;
  wire FA_out_3360;
  wire FA_out_3361;
  wire FA_out_3362;
  wire FA_out_3363;
  wire FA_out_3364;
  wire FA_out_3365;
  wire FA_out_3366;
  wire FA_out_3367;
  wire FA_out_3368;
  wire FA_out_3369;
  wire FA_out_3370;
  wire FA_out_3371;
  wire FA_out_3372;
  wire FA_out_3373;
  wire FA_out_3374;
  wire FA_out_3375;
  wire FA_out_3376;
  wire FA_out_3377;
  wire FA_out_3378;
  wire FA_out_3379;
  wire FA_out_3380;
  wire FA_out_3381;
  wire FA_out_3382;
  wire FA_out_3383;
  wire FA_out_3384;
  wire FA_out_3385;
  wire FA_out_3386;
  wire FA_out_3387;
  wire FA_out_3388;
  wire FA_out_3389;
  wire FA_out_3390;
  wire FA_out_3391;
  wire FA_out_3392;
  wire FA_out_3393;
  wire FA_out_3394;
  wire FA_out_3395;
  wire FA_out_3396;
  wire FA_out_3397;
  wire FA_out_3398;
  wire FA_out_3399;
  wire FA_out_3400;
  wire FA_out_3401;
  wire FA_out_3402;
  wire FA_out_3403;
  wire FA_out_3404;
  wire FA_out_3405;
  wire FA_out_3406;
  wire FA_out_3407;
  wire FA_out_3408;
  wire FA_out_3409;
  wire FA_out_3410;
  wire FA_out_3411;
  wire FA_out_3412;
  wire FA_out_3413;
  wire FA_out_3414;
  wire FA_out_3415;
  wire FA_out_3416;
  wire FA_out_3417;
  wire FA_out_3418;
  wire FA_out_3419;
  wire FA_out_3420;
  wire FA_out_3421;
  wire FA_out_3422;
  wire FA_out_3423;
  wire FA_out_3424;
  wire FA_out_3425;
  wire FA_out_3426;
  wire FA_out_3427;
  wire FA_out_3428;
  wire FA_out_3429;
  wire FA_out_3430;
  wire FA_out_3431;
  wire FA_out_3432;
  wire FA_out_3433;
  wire FA_out_3434;
  wire FA_out_3435;
  wire FA_out_3436;
  wire FA_out_3437;
  wire FA_out_3438;
  wire FA_out_3439;
  wire FA_out_3440;
  wire FA_out_3441;
  wire FA_out_3442;
  wire FA_out_3443;
  wire FA_out_3444;
  wire FA_out_3445;
  wire FA_out_3446;
  wire FA_out_3447;
  wire FA_out_3448;
  wire FA_out_3449;
  wire FA_out_3450;
  wire FA_out_3451;
  wire FA_out_3452;
  wire FA_out_3453;
  wire FA_out_3454;
  wire FA_out_3455;
  wire FA_out_3456;
  wire FA_out_3457;
  wire FA_out_3458;
  wire FA_out_3459;
  wire FA_out_3460;
  wire FA_out_3461;
  wire FA_out_3462;
  wire FA_out_3463;
  wire FA_out_3464;
  wire FA_out_3465;
  wire FA_out_3466;
  wire FA_out_3467;
  wire FA_out_3468;
  wire FA_out_3469;
  wire FA_out_3470;
  wire FA_out_3471;
  wire FA_out_3472;
  wire FA_out_3473;
  wire FA_out_3474;
  wire FA_out_3475;
  wire FA_out_3476;
  wire FA_out_3477;
  wire FA_out_3478;
  wire FA_out_3479;
  wire FA_out_3480;
  wire FA_out_3481;
  wire FA_out_3482;
  wire FA_out_3483;
  wire FA_out_3484;
  wire FA_out_3485;
  wire FA_out_3486;
  wire FA_out_3487;
  wire FA_out_3488;
  wire FA_out_3489;
  wire FA_out_3490;
  wire FA_out_3491;
  wire FA_out_3492;
  wire FA_out_3493;
  wire FA_out_3494;
  wire FA_out_3495;
  wire FA_out_3496;
  wire FA_out_3497;
  wire FA_out_3498;
  wire FA_out_3499;
  wire FA_out_3500;
  wire FA_out_3501;
  wire FA_out_3502;
  wire FA_out_3503;
  wire FA_out_3504;
  wire FA_out_3505;
  wire FA_out_3506;
  wire FA_out_3507;
  wire FA_out_3508;
  wire FA_out_3509;
  wire FA_out_3510;
  wire FA_out_3511;
  wire FA_out_3512;
  wire FA_out_3513;
  wire FA_out_3514;
  wire FA_out_3515;
  wire FA_out_3516;
  wire FA_out_3517;
  wire FA_out_3518;
  wire FA_out_3519;
  wire FA_out_3520;
  wire FA_out_3521;
  wire FA_out_3522;
  wire FA_out_3523;
  wire FA_out_3524;
  wire FA_out_3525;
  wire FA_out_3526;
  wire FA_out_3527;
  wire FA_out_3528;
  wire FA_out_3529;
  wire FA_out_3530;
  wire FA_out_3531;
  wire FA_out_3532;
  wire FA_out_3533;
  wire FA_out_3534;
  wire FA_out_3535;
  wire FA_out_3536;
  wire FA_out_3537;
  wire FA_out_3538;
  wire FA_out_3539;
  wire FA_out_3540;
  wire FA_out_3541;
  wire FA_out_3542;
  wire FA_out_3543;
  wire FA_out_3544;
  wire FA_out_3545;
  wire FA_out_3546;
  wire FA_out_3547;
  wire FA_out_3548;
  wire FA_out_3549;
  wire FA_out_3550;
  wire FA_out_3551;
  wire FA_out_3552;
  wire FA_out_3553;
  wire FA_out_3554;
  wire FA_out_3555;
  wire FA_out_3556;
  wire FA_out_3557;
  wire FA_out_3558;
  wire FA_out_3559;
  wire FA_out_3560;
  wire FA_out_3561;
  wire FA_out_3562;
  wire FA_out_3563;
  wire FA_out_3564;
  wire FA_out_3565;
  wire FA_out_3566;
  wire FA_out_3567;
  wire FA_out_3568;
  wire FA_out_3569;
  wire FA_out_3570;
  wire FA_out_3571;
  wire FA_out_3572;
  wire FA_out_3573;
  wire FA_out_3574;
  wire FA_out_3575;
  wire FA_out_3576;
  wire FA_out_3577;
  wire FA_out_3578;
  wire FA_out_3579;
  wire FA_out_3580;
  wire FA_out_3581;
  wire FA_out_3582;
  wire FA_out_3583;
  wire FA_out_3584;
  wire FA_out_3585;
  wire FA_out_3586;
  wire FA_out_3587;
  wire FA_out_3588;
  wire FA_out_3589;
  wire FA_out_3590;
  wire FA_out_3591;
  wire FA_out_3592;
  wire FA_out_3593;
  wire FA_out_3594;
  wire FA_out_3595;
  wire FA_out_3596;
  wire FA_out_3597;
  wire FA_out_3598;
  wire FA_out_3599;
  wire FA_out_3600;
  wire FA_out_3601;
  wire FA_out_3602;
  wire FA_out_3603;
  wire FA_out_3604;
  wire FA_out_3605;
  wire FA_out_3606;
  wire FA_out_3607;
  wire FA_out_3608;
  wire FA_out_3609;
  wire FA_out_3610;
  wire FA_out_3611;
  wire FA_out_3612;
  wire FA_out_3613;
  wire FA_out_3614;
  wire FA_out_3615;
  wire FA_out_3616;
  wire FA_out_3617;
  wire FA_out_3618;
  wire FA_out_3619;
  wire FA_out_3620;
  wire FA_out_3621;
  wire FA_out_3622;
  wire FA_out_3623;
  wire FA_out_3624;
  wire FA_out_3625;
  wire FA_out_3626;
  wire FA_out_3627;
  wire FA_out_3628;
  wire FA_out_3629;
  wire FA_out_3630;
  wire FA_out_3631;
  wire FA_out_3632;
  wire FA_out_3633;
  wire FA_out_3634;
  wire FA_out_3635;
  wire FA_out_3636;
  wire FA_out_3637;
  wire FA_out_3638;
  wire FA_out_3639;
  wire FA_out_3640;
  wire FA_out_3641;
  wire FA_out_3642;
  wire FA_out_3643;
  wire FA_out_3644;
  wire FA_out_3645;
  wire FA_out_3646;
  wire FA_out_3647;
  wire FA_out_3648;
  wire FA_out_3649;
  wire FA_out_3650;
  wire FA_out_3651;
  wire FA_out_3652;
  wire FA_out_3653;
  wire FA_out_3654;
  wire FA_out_3655;
  wire FA_out_3656;
  wire FA_out_3657;
  wire FA_out_3658;
  wire FA_out_3659;
  wire FA_out_3660;
  wire FA_out_3661;
  wire FA_out_3662;
  wire FA_out_3663;
  wire FA_out_3664;
  wire FA_out_3665;
  wire FA_out_3666;
  wire FA_out_3667;
  wire FA_out_3668;
  wire FA_out_3669;
  wire FA_out_3670;
  wire FA_out_3671;
  wire FA_out_3672;
  wire FA_out_3673;
  wire FA_out_3674;
  wire FA_out_3675;
  wire FA_out_3676;
  wire FA_out_3677;
  wire FA_out_3678;
  wire FA_out_3679;
  wire FA_out_3680;
  wire FA_out_3681;
  wire FA_out_3682;
  wire FA_out_3683;
  wire FA_out_3684;
  wire FA_out_3685;
  wire FA_out_3686;
  wire FA_out_3687;
  wire FA_out_3688;
  wire FA_out_3689;
  wire FA_out_3690;
  wire FA_out_3691;
  wire FA_out_3692;
  wire FA_out_3693;
  wire FA_out_3694;
  wire FA_out_3695;
  wire FA_out_3696;
  wire FA_out_3697;
  wire FA_out_3698;
  wire FA_out_3699;
  wire FA_out_3700;
  wire FA_out_3701;
  wire FA_out_3702;
  wire FA_out_3703;
  wire FA_out_3704;
  wire FA_out_3705;
  wire FA_out_3706;
  wire FA_out_3707;
  wire FA_out_3708;
  wire FA_out_3709;
  wire FA_out_3710;
  wire FA_out_3711;
  wire FA_out_3712;
  wire FA_out_3713;
  wire FA_out_3714;
  wire FA_out_3715;
  wire FA_out_3716;
  wire FA_out_3717;
  wire FA_out_3718;
  wire FA_out_3719;
  wire FA_out_3720;
  wire FA_out_3721;
  wire FA_out_3722;
  wire FA_out_3723;
  wire FA_out_3724;
  wire FA_out_3725;
  wire FA_out_3726;
  wire FA_out_3727;
  wire FA_out_3728;
  wire FA_out_3729;
  wire FA_out_3730;
  wire FA_out_3731;
  wire FA_out_3732;
  wire FA_out_3733;
  wire FA_out_3734;
  wire FA_out_3735;
  wire FA_out_3736;
  wire FA_out_3737;
  wire FA_out_3738;
  wire FA_out_3739;
  wire FA_out_3740;
  wire FA_out_3741;
  wire FA_out_3742;
  wire FA_out_3743;
  wire FA_out_3744;
  wire FA_out_3745;
  wire FA_out_3746;
  wire FA_out_3747;
  wire FA_out_3748;
  wire FA_out_3749;
  wire FA_out_3750;
  wire FA_out_3751;
  wire FA_out_3752;
  wire FA_out_3753;
  wire FA_out_3754;
  wire FA_out_3755;
  wire FA_out_3756;
  wire FA_out_3757;
  wire FA_out_3758;
  wire FA_out_3759;
  wire FA_out_3760;
  wire FA_out_3761;
  wire FA_out_3762;
  wire FA_out_3763;
  wire FA_out_3764;
  wire FA_out_3765;
  wire FA_out_3766;
  wire FA_out_3767;
  wire FA_out_3768;
  wire FA_out_3769;
  wire FA_out_3770;
  wire FA_out_3771;
  wire FA_out_3772;
  wire FA_out_3773;
  wire FA_out_3774;
  wire FA_out_3775;
  wire FA_out_3776;
  wire FA_out_3777;
  wire FA_out_3778;
  wire FA_out_3779;
  wire FA_out_3780;
  wire FA_out_3781;
  wire FA_out_3782;
  wire FA_out_3783;
  wire FA_out_3784;
  wire FA_out_3785;
  wire FA_out_3786;
  wire FA_out_3787;
  wire FA_out_3788;
  wire FA_out_3789;
  wire FA_out_3790;
  wire FA_out_3791;
  wire FA_out_3792;
  wire FA_out_3793;
  wire FA_out_3794;
  wire FA_out_3795;
  wire FA_out_3796;
  wire FA_out_3797;
  wire FA_out_3798;
  wire FA_out_3799;
  wire FA_out_3800;
  wire FA_out_3801;
  wire FA_out_3802;
  wire FA_out_3803;
  wire FA_out_3804;
  wire FA_out_3805;
  wire FA_out_3806;
  wire FA_out_3807;
  wire FA_out_3808;
  wire FA_out_3809;
  wire FA_out_3810;
  wire FA_out_3811;
  wire FA_out_3812;
  wire FA_out_3813;
  wire FA_out_3814;
  wire FA_out_3815;
  wire FA_out_3816;
  wire FA_out_3817;
  wire FA_out_3818;
  wire FA_out_3819;
  wire FA_out_3820;
  wire FA_out_3821;
  wire FA_out_3822;
  wire FA_out_3823;
  wire FA_out_3824;
  wire FA_out_3825;
  wire FA_out_3826;
  wire FA_out_3827;
  wire FA_out_3828;
  wire FA_out_3829;
  wire FA_out_3830;
  wire FA_out_3831;
  wire FA_out_3832;
  wire FA_out_3833;
  wire FA_out_3834;
  wire FA_out_3835;
  wire FA_out_3836;
  wire FA_out_3837;
  wire FA_out_3838;
  wire FA_out_3839;
  wire FA_out_3840;
  wire FA_out_3841;
  wire FA_out_3842;
  wire FA_out_3843;
  wire FA_cout_0;
  wire FA_cout_1;
  wire FA_cout_2;
  wire FA_cout_3;
  wire FA_cout_4;
  wire FA_cout_5;
  wire FA_cout_6;
  wire FA_cout_7;
  wire FA_cout_8;
  wire FA_cout_9;
  wire FA_cout_10;
  wire FA_cout_11;
  wire FA_cout_12;
  wire FA_cout_13;
  wire FA_cout_14;
  wire FA_cout_15;
  wire FA_cout_16;
  wire FA_cout_17;
  wire FA_cout_18;
  wire FA_cout_19;
  wire FA_cout_20;
  wire FA_cout_21;
  wire FA_cout_22;
  wire FA_cout_23;
  wire FA_cout_24;
  wire FA_cout_25;
  wire FA_cout_26;
  wire FA_cout_27;
  wire FA_cout_28;
  wire FA_cout_29;
  wire FA_cout_30;
  wire FA_cout_31;
  wire FA_cout_32;
  wire FA_cout_33;
  wire FA_cout_34;
  wire FA_cout_35;
  wire FA_cout_36;
  wire FA_cout_37;
  wire FA_cout_38;
  wire FA_cout_39;
  wire FA_cout_40;
  wire FA_cout_41;
  wire FA_cout_42;
  wire FA_cout_43;
  wire FA_cout_44;
  wire FA_cout_45;
  wire FA_cout_46;
  wire FA_cout_47;
  wire FA_cout_48;
  wire FA_cout_49;
  wire FA_cout_50;
  wire FA_cout_51;
  wire FA_cout_52;
  wire FA_cout_53;
  wire FA_cout_54;
  wire FA_cout_55;
  wire FA_cout_56;
  wire FA_cout_57;
  wire FA_cout_58;
  wire FA_cout_59;
  wire FA_cout_60;
  wire FA_cout_61;
  wire FA_cout_62;
  wire FA_cout_63;
  wire FA_cout_64;
  wire FA_cout_65;
  wire FA_cout_66;
  wire FA_cout_67;
  wire FA_cout_68;
  wire FA_cout_69;
  wire FA_cout_70;
  wire FA_cout_71;
  wire FA_cout_72;
  wire FA_cout_73;
  wire FA_cout_74;
  wire FA_cout_75;
  wire FA_cout_76;
  wire FA_cout_77;
  wire FA_cout_78;
  wire FA_cout_79;
  wire FA_cout_80;
  wire FA_cout_81;
  wire FA_cout_82;
  wire FA_cout_83;
  wire FA_cout_84;
  wire FA_cout_85;
  wire FA_cout_86;
  wire FA_cout_87;
  wire FA_cout_88;
  wire FA_cout_89;
  wire FA_cout_90;
  wire FA_cout_91;
  wire FA_cout_92;
  wire FA_cout_93;
  wire FA_cout_94;
  wire FA_cout_95;
  wire FA_cout_96;
  wire FA_cout_97;
  wire FA_cout_98;
  wire FA_cout_99;
  wire FA_cout_100;
  wire FA_cout_101;
  wire FA_cout_102;
  wire FA_cout_103;
  wire FA_cout_104;
  wire FA_cout_105;
  wire FA_cout_106;
  wire FA_cout_107;
  wire FA_cout_108;
  wire FA_cout_109;
  wire FA_cout_110;
  wire FA_cout_111;
  wire FA_cout_112;
  wire FA_cout_113;
  wire FA_cout_114;
  wire FA_cout_115;
  wire FA_cout_116;
  wire FA_cout_117;
  wire FA_cout_118;
  wire FA_cout_119;
  wire FA_cout_120;
  wire FA_cout_121;
  wire FA_cout_122;
  wire FA_cout_123;
  wire FA_cout_124;
  wire FA_cout_125;
  wire FA_cout_126;
  wire FA_cout_127;
  wire FA_cout_128;
  wire FA_cout_129;
  wire FA_cout_130;
  wire FA_cout_131;
  wire FA_cout_132;
  wire FA_cout_133;
  wire FA_cout_134;
  wire FA_cout_135;
  wire FA_cout_136;
  wire FA_cout_137;
  wire FA_cout_138;
  wire FA_cout_139;
  wire FA_cout_140;
  wire FA_cout_141;
  wire FA_cout_142;
  wire FA_cout_143;
  wire FA_cout_144;
  wire FA_cout_145;
  wire FA_cout_146;
  wire FA_cout_147;
  wire FA_cout_148;
  wire FA_cout_149;
  wire FA_cout_150;
  wire FA_cout_151;
  wire FA_cout_152;
  wire FA_cout_153;
  wire FA_cout_154;
  wire FA_cout_155;
  wire FA_cout_156;
  wire FA_cout_157;
  wire FA_cout_158;
  wire FA_cout_159;
  wire FA_cout_160;
  wire FA_cout_161;
  wire FA_cout_162;
  wire FA_cout_163;
  wire FA_cout_164;
  wire FA_cout_165;
  wire FA_cout_166;
  wire FA_cout_167;
  wire FA_cout_168;
  wire FA_cout_169;
  wire FA_cout_170;
  wire FA_cout_171;
  wire FA_cout_172;
  wire FA_cout_173;
  wire FA_cout_174;
  wire FA_cout_175;
  wire FA_cout_176;
  wire FA_cout_177;
  wire FA_cout_178;
  wire FA_cout_179;
  wire FA_cout_180;
  wire FA_cout_181;
  wire FA_cout_182;
  wire FA_cout_183;
  wire FA_cout_184;
  wire FA_cout_185;
  wire FA_cout_186;
  wire FA_cout_187;
  wire FA_cout_188;
  wire FA_cout_189;
  wire FA_cout_190;
  wire FA_cout_191;
  wire FA_cout_192;
  wire FA_cout_193;
  wire FA_cout_194;
  wire FA_cout_195;
  wire FA_cout_196;
  wire FA_cout_197;
  wire FA_cout_198;
  wire FA_cout_199;
  wire FA_cout_200;
  wire FA_cout_201;
  wire FA_cout_202;
  wire FA_cout_203;
  wire FA_cout_204;
  wire FA_cout_205;
  wire FA_cout_206;
  wire FA_cout_207;
  wire FA_cout_208;
  wire FA_cout_209;
  wire FA_cout_210;
  wire FA_cout_211;
  wire FA_cout_212;
  wire FA_cout_213;
  wire FA_cout_214;
  wire FA_cout_215;
  wire FA_cout_216;
  wire FA_cout_217;
  wire FA_cout_218;
  wire FA_cout_219;
  wire FA_cout_220;
  wire FA_cout_221;
  wire FA_cout_222;
  wire FA_cout_223;
  wire FA_cout_224;
  wire FA_cout_225;
  wire FA_cout_226;
  wire FA_cout_227;
  wire FA_cout_228;
  wire FA_cout_229;
  wire FA_cout_230;
  wire FA_cout_231;
  wire FA_cout_232;
  wire FA_cout_233;
  wire FA_cout_234;
  wire FA_cout_235;
  wire FA_cout_236;
  wire FA_cout_237;
  wire FA_cout_238;
  wire FA_cout_239;
  wire FA_cout_240;
  wire FA_cout_241;
  wire FA_cout_242;
  wire FA_cout_243;
  wire FA_cout_244;
  wire FA_cout_245;
  wire FA_cout_246;
  wire FA_cout_247;
  wire FA_cout_248;
  wire FA_cout_249;
  wire FA_cout_250;
  wire FA_cout_251;
  wire FA_cout_252;
  wire FA_cout_253;
  wire FA_cout_254;
  wire FA_cout_255;
  wire FA_cout_256;
  wire FA_cout_257;
  wire FA_cout_258;
  wire FA_cout_259;
  wire FA_cout_260;
  wire FA_cout_261;
  wire FA_cout_262;
  wire FA_cout_263;
  wire FA_cout_264;
  wire FA_cout_265;
  wire FA_cout_266;
  wire FA_cout_267;
  wire FA_cout_268;
  wire FA_cout_269;
  wire FA_cout_270;
  wire FA_cout_271;
  wire FA_cout_272;
  wire FA_cout_273;
  wire FA_cout_274;
  wire FA_cout_275;
  wire FA_cout_276;
  wire FA_cout_277;
  wire FA_cout_278;
  wire FA_cout_279;
  wire FA_cout_280;
  wire FA_cout_281;
  wire FA_cout_282;
  wire FA_cout_283;
  wire FA_cout_284;
  wire FA_cout_285;
  wire FA_cout_286;
  wire FA_cout_287;
  wire FA_cout_288;
  wire FA_cout_289;
  wire FA_cout_290;
  wire FA_cout_291;
  wire FA_cout_292;
  wire FA_cout_293;
  wire FA_cout_294;
  wire FA_cout_295;
  wire FA_cout_296;
  wire FA_cout_297;
  wire FA_cout_298;
  wire FA_cout_299;
  wire FA_cout_300;
  wire FA_cout_301;
  wire FA_cout_302;
  wire FA_cout_303;
  wire FA_cout_304;
  wire FA_cout_305;
  wire FA_cout_306;
  wire FA_cout_307;
  wire FA_cout_308;
  wire FA_cout_309;
  wire FA_cout_310;
  wire FA_cout_311;
  wire FA_cout_312;
  wire FA_cout_313;
  wire FA_cout_314;
  wire FA_cout_315;
  wire FA_cout_316;
  wire FA_cout_317;
  wire FA_cout_318;
  wire FA_cout_319;
  wire FA_cout_320;
  wire FA_cout_321;
  wire FA_cout_322;
  wire FA_cout_323;
  wire FA_cout_324;
  wire FA_cout_325;
  wire FA_cout_326;
  wire FA_cout_327;
  wire FA_cout_328;
  wire FA_cout_329;
  wire FA_cout_330;
  wire FA_cout_331;
  wire FA_cout_332;
  wire FA_cout_333;
  wire FA_cout_334;
  wire FA_cout_335;
  wire FA_cout_336;
  wire FA_cout_337;
  wire FA_cout_338;
  wire FA_cout_339;
  wire FA_cout_340;
  wire FA_cout_341;
  wire FA_cout_342;
  wire FA_cout_343;
  wire FA_cout_344;
  wire FA_cout_345;
  wire FA_cout_346;
  wire FA_cout_347;
  wire FA_cout_348;
  wire FA_cout_349;
  wire FA_cout_350;
  wire FA_cout_351;
  wire FA_cout_352;
  wire FA_cout_353;
  wire FA_cout_354;
  wire FA_cout_355;
  wire FA_cout_356;
  wire FA_cout_357;
  wire FA_cout_358;
  wire FA_cout_359;
  wire FA_cout_360;
  wire FA_cout_361;
  wire FA_cout_362;
  wire FA_cout_363;
  wire FA_cout_364;
  wire FA_cout_365;
  wire FA_cout_366;
  wire FA_cout_367;
  wire FA_cout_368;
  wire FA_cout_369;
  wire FA_cout_370;
  wire FA_cout_371;
  wire FA_cout_372;
  wire FA_cout_373;
  wire FA_cout_374;
  wire FA_cout_375;
  wire FA_cout_376;
  wire FA_cout_377;
  wire FA_cout_378;
  wire FA_cout_379;
  wire FA_cout_380;
  wire FA_cout_381;
  wire FA_cout_382;
  wire FA_cout_383;
  wire FA_cout_384;
  wire FA_cout_385;
  wire FA_cout_386;
  wire FA_cout_387;
  wire FA_cout_388;
  wire FA_cout_389;
  wire FA_cout_390;
  wire FA_cout_391;
  wire FA_cout_392;
  wire FA_cout_393;
  wire FA_cout_394;
  wire FA_cout_395;
  wire FA_cout_396;
  wire FA_cout_397;
  wire FA_cout_398;
  wire FA_cout_399;
  wire FA_cout_400;
  wire FA_cout_401;
  wire FA_cout_402;
  wire FA_cout_403;
  wire FA_cout_404;
  wire FA_cout_405;
  wire FA_cout_406;
  wire FA_cout_407;
  wire FA_cout_408;
  wire FA_cout_409;
  wire FA_cout_410;
  wire FA_cout_411;
  wire FA_cout_412;
  wire FA_cout_413;
  wire FA_cout_414;
  wire FA_cout_415;
  wire FA_cout_416;
  wire FA_cout_417;
  wire FA_cout_418;
  wire FA_cout_419;
  wire FA_cout_420;
  wire FA_cout_421;
  wire FA_cout_422;
  wire FA_cout_423;
  wire FA_cout_424;
  wire FA_cout_425;
  wire FA_cout_426;
  wire FA_cout_427;
  wire FA_cout_428;
  wire FA_cout_429;
  wire FA_cout_430;
  wire FA_cout_431;
  wire FA_cout_432;
  wire FA_cout_433;
  wire FA_cout_434;
  wire FA_cout_435;
  wire FA_cout_436;
  wire FA_cout_437;
  wire FA_cout_438;
  wire FA_cout_439;
  wire FA_cout_440;
  wire FA_cout_441;
  wire FA_cout_442;
  wire FA_cout_443;
  wire FA_cout_444;
  wire FA_cout_445;
  wire FA_cout_446;
  wire FA_cout_447;
  wire FA_cout_448;
  wire FA_cout_449;
  wire FA_cout_450;
  wire FA_cout_451;
  wire FA_cout_452;
  wire FA_cout_453;
  wire FA_cout_454;
  wire FA_cout_455;
  wire FA_cout_456;
  wire FA_cout_457;
  wire FA_cout_458;
  wire FA_cout_459;
  wire FA_cout_460;
  wire FA_cout_461;
  wire FA_cout_462;
  wire FA_cout_463;
  wire FA_cout_464;
  wire FA_cout_465;
  wire FA_cout_466;
  wire FA_cout_467;
  wire FA_cout_468;
  wire FA_cout_469;
  wire FA_cout_470;
  wire FA_cout_471;
  wire FA_cout_472;
  wire FA_cout_473;
  wire FA_cout_474;
  wire FA_cout_475;
  wire FA_cout_476;
  wire FA_cout_477;
  wire FA_cout_478;
  wire FA_cout_479;
  wire FA_cout_480;
  wire FA_cout_481;
  wire FA_cout_482;
  wire FA_cout_483;
  wire FA_cout_484;
  wire FA_cout_485;
  wire FA_cout_486;
  wire FA_cout_487;
  wire FA_cout_488;
  wire FA_cout_489;
  wire FA_cout_490;
  wire FA_cout_491;
  wire FA_cout_492;
  wire FA_cout_493;
  wire FA_cout_494;
  wire FA_cout_495;
  wire FA_cout_496;
  wire FA_cout_497;
  wire FA_cout_498;
  wire FA_cout_499;
  wire FA_cout_500;
  wire FA_cout_501;
  wire FA_cout_502;
  wire FA_cout_503;
  wire FA_cout_504;
  wire FA_cout_505;
  wire FA_cout_506;
  wire FA_cout_507;
  wire FA_cout_508;
  wire FA_cout_509;
  wire FA_cout_510;
  wire FA_cout_511;
  wire FA_cout_512;
  wire FA_cout_513;
  wire FA_cout_514;
  wire FA_cout_515;
  wire FA_cout_516;
  wire FA_cout_517;
  wire FA_cout_518;
  wire FA_cout_519;
  wire FA_cout_520;
  wire FA_cout_521;
  wire FA_cout_522;
  wire FA_cout_523;
  wire FA_cout_524;
  wire FA_cout_525;
  wire FA_cout_526;
  wire FA_cout_527;
  wire FA_cout_528;
  wire FA_cout_529;
  wire FA_cout_530;
  wire FA_cout_531;
  wire FA_cout_532;
  wire FA_cout_533;
  wire FA_cout_534;
  wire FA_cout_535;
  wire FA_cout_536;
  wire FA_cout_537;
  wire FA_cout_538;
  wire FA_cout_539;
  wire FA_cout_540;
  wire FA_cout_541;
  wire FA_cout_542;
  wire FA_cout_543;
  wire FA_cout_544;
  wire FA_cout_545;
  wire FA_cout_546;
  wire FA_cout_547;
  wire FA_cout_548;
  wire FA_cout_549;
  wire FA_cout_550;
  wire FA_cout_551;
  wire FA_cout_552;
  wire FA_cout_553;
  wire FA_cout_554;
  wire FA_cout_555;
  wire FA_cout_556;
  wire FA_cout_557;
  wire FA_cout_558;
  wire FA_cout_559;
  wire FA_cout_560;
  wire FA_cout_561;
  wire FA_cout_562;
  wire FA_cout_563;
  wire FA_cout_564;
  wire FA_cout_565;
  wire FA_cout_566;
  wire FA_cout_567;
  wire FA_cout_568;
  wire FA_cout_569;
  wire FA_cout_570;
  wire FA_cout_571;
  wire FA_cout_572;
  wire FA_cout_573;
  wire FA_cout_574;
  wire FA_cout_575;
  wire FA_cout_576;
  wire FA_cout_577;
  wire FA_cout_578;
  wire FA_cout_579;
  wire FA_cout_580;
  wire FA_cout_581;
  wire FA_cout_582;
  wire FA_cout_583;
  wire FA_cout_584;
  wire FA_cout_585;
  wire FA_cout_586;
  wire FA_cout_587;
  wire FA_cout_588;
  wire FA_cout_589;
  wire FA_cout_590;
  wire FA_cout_591;
  wire FA_cout_592;
  wire FA_cout_593;
  wire FA_cout_594;
  wire FA_cout_595;
  wire FA_cout_596;
  wire FA_cout_597;
  wire FA_cout_598;
  wire FA_cout_599;
  wire FA_cout_600;
  wire FA_cout_601;
  wire FA_cout_602;
  wire FA_cout_603;
  wire FA_cout_604;
  wire FA_cout_605;
  wire FA_cout_606;
  wire FA_cout_607;
  wire FA_cout_608;
  wire FA_cout_609;
  wire FA_cout_610;
  wire FA_cout_611;
  wire FA_cout_612;
  wire FA_cout_613;
  wire FA_cout_614;
  wire FA_cout_615;
  wire FA_cout_616;
  wire FA_cout_617;
  wire FA_cout_618;
  wire FA_cout_619;
  wire FA_cout_620;
  wire FA_cout_621;
  wire FA_cout_622;
  wire FA_cout_623;
  wire FA_cout_624;
  wire FA_cout_625;
  wire FA_cout_626;
  wire FA_cout_627;
  wire FA_cout_628;
  wire FA_cout_629;
  wire FA_cout_630;
  wire FA_cout_631;
  wire FA_cout_632;
  wire FA_cout_633;
  wire FA_cout_634;
  wire FA_cout_635;
  wire FA_cout_636;
  wire FA_cout_637;
  wire FA_cout_638;
  wire FA_cout_639;
  wire FA_cout_640;
  wire FA_cout_641;
  wire FA_cout_642;
  wire FA_cout_643;
  wire FA_cout_644;
  wire FA_cout_645;
  wire FA_cout_646;
  wire FA_cout_647;
  wire FA_cout_648;
  wire FA_cout_649;
  wire FA_cout_650;
  wire FA_cout_651;
  wire FA_cout_652;
  wire FA_cout_653;
  wire FA_cout_654;
  wire FA_cout_655;
  wire FA_cout_656;
  wire FA_cout_657;
  wire FA_cout_658;
  wire FA_cout_659;
  wire FA_cout_660;
  wire FA_cout_661;
  wire FA_cout_662;
  wire FA_cout_663;
  wire FA_cout_664;
  wire FA_cout_665;
  wire FA_cout_666;
  wire FA_cout_667;
  wire FA_cout_668;
  wire FA_cout_669;
  wire FA_cout_670;
  wire FA_cout_671;
  wire FA_cout_672;
  wire FA_cout_673;
  wire FA_cout_674;
  wire FA_cout_675;
  wire FA_cout_676;
  wire FA_cout_677;
  wire FA_cout_678;
  wire FA_cout_679;
  wire FA_cout_680;
  wire FA_cout_681;
  wire FA_cout_682;
  wire FA_cout_683;
  wire FA_cout_684;
  wire FA_cout_685;
  wire FA_cout_686;
  wire FA_cout_687;
  wire FA_cout_688;
  wire FA_cout_689;
  wire FA_cout_690;
  wire FA_cout_691;
  wire FA_cout_692;
  wire FA_cout_693;
  wire FA_cout_694;
  wire FA_cout_695;
  wire FA_cout_696;
  wire FA_cout_697;
  wire FA_cout_698;
  wire FA_cout_699;
  wire FA_cout_700;
  wire FA_cout_701;
  wire FA_cout_702;
  wire FA_cout_703;
  wire FA_cout_704;
  wire FA_cout_705;
  wire FA_cout_706;
  wire FA_cout_707;
  wire FA_cout_708;
  wire FA_cout_709;
  wire FA_cout_710;
  wire FA_cout_711;
  wire FA_cout_712;
  wire FA_cout_713;
  wire FA_cout_714;
  wire FA_cout_715;
  wire FA_cout_716;
  wire FA_cout_717;
  wire FA_cout_718;
  wire FA_cout_719;
  wire FA_cout_720;
  wire FA_cout_721;
  wire FA_cout_722;
  wire FA_cout_723;
  wire FA_cout_724;
  wire FA_cout_725;
  wire FA_cout_726;
  wire FA_cout_727;
  wire FA_cout_728;
  wire FA_cout_729;
  wire FA_cout_730;
  wire FA_cout_731;
  wire FA_cout_732;
  wire FA_cout_733;
  wire FA_cout_734;
  wire FA_cout_735;
  wire FA_cout_736;
  wire FA_cout_737;
  wire FA_cout_738;
  wire FA_cout_739;
  wire FA_cout_740;
  wire FA_cout_741;
  wire FA_cout_742;
  wire FA_cout_743;
  wire FA_cout_744;
  wire FA_cout_745;
  wire FA_cout_746;
  wire FA_cout_747;
  wire FA_cout_748;
  wire FA_cout_749;
  wire FA_cout_750;
  wire FA_cout_751;
  wire FA_cout_752;
  wire FA_cout_753;
  wire FA_cout_754;
  wire FA_cout_755;
  wire FA_cout_756;
  wire FA_cout_757;
  wire FA_cout_758;
  wire FA_cout_759;
  wire FA_cout_760;
  wire FA_cout_761;
  wire FA_cout_762;
  wire FA_cout_763;
  wire FA_cout_764;
  wire FA_cout_765;
  wire FA_cout_766;
  wire FA_cout_767;
  wire FA_cout_768;
  wire FA_cout_769;
  wire FA_cout_770;
  wire FA_cout_771;
  wire FA_cout_772;
  wire FA_cout_773;
  wire FA_cout_774;
  wire FA_cout_775;
  wire FA_cout_776;
  wire FA_cout_777;
  wire FA_cout_778;
  wire FA_cout_779;
  wire FA_cout_780;
  wire FA_cout_781;
  wire FA_cout_782;
  wire FA_cout_783;
  wire FA_cout_784;
  wire FA_cout_785;
  wire FA_cout_786;
  wire FA_cout_787;
  wire FA_cout_788;
  wire FA_cout_789;
  wire FA_cout_790;
  wire FA_cout_791;
  wire FA_cout_792;
  wire FA_cout_793;
  wire FA_cout_794;
  wire FA_cout_795;
  wire FA_cout_796;
  wire FA_cout_797;
  wire FA_cout_798;
  wire FA_cout_799;
  wire FA_cout_800;
  wire FA_cout_801;
  wire FA_cout_802;
  wire FA_cout_803;
  wire FA_cout_804;
  wire FA_cout_805;
  wire FA_cout_806;
  wire FA_cout_807;
  wire FA_cout_808;
  wire FA_cout_809;
  wire FA_cout_810;
  wire FA_cout_811;
  wire FA_cout_812;
  wire FA_cout_813;
  wire FA_cout_814;
  wire FA_cout_815;
  wire FA_cout_816;
  wire FA_cout_817;
  wire FA_cout_818;
  wire FA_cout_819;
  wire FA_cout_820;
  wire FA_cout_821;
  wire FA_cout_822;
  wire FA_cout_823;
  wire FA_cout_824;
  wire FA_cout_825;
  wire FA_cout_826;
  wire FA_cout_827;
  wire FA_cout_828;
  wire FA_cout_829;
  wire FA_cout_830;
  wire FA_cout_831;
  wire FA_cout_832;
  wire FA_cout_833;
  wire FA_cout_834;
  wire FA_cout_835;
  wire FA_cout_836;
  wire FA_cout_837;
  wire FA_cout_838;
  wire FA_cout_839;
  wire FA_cout_840;
  wire FA_cout_841;
  wire FA_cout_842;
  wire FA_cout_843;
  wire FA_cout_844;
  wire FA_cout_845;
  wire FA_cout_846;
  wire FA_cout_847;
  wire FA_cout_848;
  wire FA_cout_849;
  wire FA_cout_850;
  wire FA_cout_851;
  wire FA_cout_852;
  wire FA_cout_853;
  wire FA_cout_854;
  wire FA_cout_855;
  wire FA_cout_856;
  wire FA_cout_857;
  wire FA_cout_858;
  wire FA_cout_859;
  wire FA_cout_860;
  wire FA_cout_861;
  wire FA_cout_862;
  wire FA_cout_863;
  wire FA_cout_864;
  wire FA_cout_865;
  wire FA_cout_866;
  wire FA_cout_867;
  wire FA_cout_868;
  wire FA_cout_869;
  wire FA_cout_870;
  wire FA_cout_871;
  wire FA_cout_872;
  wire FA_cout_873;
  wire FA_cout_874;
  wire FA_cout_875;
  wire FA_cout_876;
  wire FA_cout_877;
  wire FA_cout_878;
  wire FA_cout_879;
  wire FA_cout_880;
  wire FA_cout_881;
  wire FA_cout_882;
  wire FA_cout_883;
  wire FA_cout_884;
  wire FA_cout_885;
  wire FA_cout_886;
  wire FA_cout_887;
  wire FA_cout_888;
  wire FA_cout_889;
  wire FA_cout_890;
  wire FA_cout_891;
  wire FA_cout_892;
  wire FA_cout_893;
  wire FA_cout_894;
  wire FA_cout_895;
  wire FA_cout_896;
  wire FA_cout_897;
  wire FA_cout_898;
  wire FA_cout_899;
  wire FA_cout_900;
  wire FA_cout_901;
  wire FA_cout_902;
  wire FA_cout_903;
  wire FA_cout_904;
  wire FA_cout_905;
  wire FA_cout_906;
  wire FA_cout_907;
  wire FA_cout_908;
  wire FA_cout_909;
  wire FA_cout_910;
  wire FA_cout_911;
  wire FA_cout_912;
  wire FA_cout_913;
  wire FA_cout_914;
  wire FA_cout_915;
  wire FA_cout_916;
  wire FA_cout_917;
  wire FA_cout_918;
  wire FA_cout_919;
  wire FA_cout_920;
  wire FA_cout_921;
  wire FA_cout_922;
  wire FA_cout_923;
  wire FA_cout_924;
  wire FA_cout_925;
  wire FA_cout_926;
  wire FA_cout_927;
  wire FA_cout_928;
  wire FA_cout_929;
  wire FA_cout_930;
  wire FA_cout_931;
  wire FA_cout_932;
  wire FA_cout_933;
  wire FA_cout_934;
  wire FA_cout_935;
  wire FA_cout_936;
  wire FA_cout_937;
  wire FA_cout_938;
  wire FA_cout_939;
  wire FA_cout_940;
  wire FA_cout_941;
  wire FA_cout_942;
  wire FA_cout_943;
  wire FA_cout_944;
  wire FA_cout_945;
  wire FA_cout_946;
  wire FA_cout_947;
  wire FA_cout_948;
  wire FA_cout_949;
  wire FA_cout_950;
  wire FA_cout_951;
  wire FA_cout_952;
  wire FA_cout_953;
  wire FA_cout_954;
  wire FA_cout_955;
  wire FA_cout_956;
  wire FA_cout_957;
  wire FA_cout_958;
  wire FA_cout_959;
  wire FA_cout_960;
  wire FA_cout_961;
  wire FA_cout_962;
  wire FA_cout_963;
  wire FA_cout_964;
  wire FA_cout_965;
  wire FA_cout_966;
  wire FA_cout_967;
  wire FA_cout_968;
  wire FA_cout_969;
  wire FA_cout_970;
  wire FA_cout_971;
  wire FA_cout_972;
  wire FA_cout_973;
  wire FA_cout_974;
  wire FA_cout_975;
  wire FA_cout_976;
  wire FA_cout_977;
  wire FA_cout_978;
  wire FA_cout_979;
  wire FA_cout_980;
  wire FA_cout_981;
  wire FA_cout_982;
  wire FA_cout_983;
  wire FA_cout_984;
  wire FA_cout_985;
  wire FA_cout_986;
  wire FA_cout_987;
  wire FA_cout_988;
  wire FA_cout_989;
  wire FA_cout_990;
  wire FA_cout_991;
  wire FA_cout_992;
  wire FA_cout_993;
  wire FA_cout_994;
  wire FA_cout_995;
  wire FA_cout_996;
  wire FA_cout_997;
  wire FA_cout_998;
  wire FA_cout_999;
  wire FA_cout_1000;
  wire FA_cout_1001;
  wire FA_cout_1002;
  wire FA_cout_1003;
  wire FA_cout_1004;
  wire FA_cout_1005;
  wire FA_cout_1006;
  wire FA_cout_1007;
  wire FA_cout_1008;
  wire FA_cout_1009;
  wire FA_cout_1010;
  wire FA_cout_1011;
  wire FA_cout_1012;
  wire FA_cout_1013;
  wire FA_cout_1014;
  wire FA_cout_1015;
  wire FA_cout_1016;
  wire FA_cout_1017;
  wire FA_cout_1018;
  wire FA_cout_1019;
  wire FA_cout_1020;
  wire FA_cout_1021;
  wire FA_cout_1022;
  wire FA_cout_1023;
  wire FA_cout_1024;
  wire FA_cout_1025;
  wire FA_cout_1026;
  wire FA_cout_1027;
  wire FA_cout_1028;
  wire FA_cout_1029;
  wire FA_cout_1030;
  wire FA_cout_1031;
  wire FA_cout_1032;
  wire FA_cout_1033;
  wire FA_cout_1034;
  wire FA_cout_1035;
  wire FA_cout_1036;
  wire FA_cout_1037;
  wire FA_cout_1038;
  wire FA_cout_1039;
  wire FA_cout_1040;
  wire FA_cout_1041;
  wire FA_cout_1042;
  wire FA_cout_1043;
  wire FA_cout_1044;
  wire FA_cout_1045;
  wire FA_cout_1046;
  wire FA_cout_1047;
  wire FA_cout_1048;
  wire FA_cout_1049;
  wire FA_cout_1050;
  wire FA_cout_1051;
  wire FA_cout_1052;
  wire FA_cout_1053;
  wire FA_cout_1054;
  wire FA_cout_1055;
  wire FA_cout_1056;
  wire FA_cout_1057;
  wire FA_cout_1058;
  wire FA_cout_1059;
  wire FA_cout_1060;
  wire FA_cout_1061;
  wire FA_cout_1062;
  wire FA_cout_1063;
  wire FA_cout_1064;
  wire FA_cout_1065;
  wire FA_cout_1066;
  wire FA_cout_1067;
  wire FA_cout_1068;
  wire FA_cout_1069;
  wire FA_cout_1070;
  wire FA_cout_1071;
  wire FA_cout_1072;
  wire FA_cout_1073;
  wire FA_cout_1074;
  wire FA_cout_1075;
  wire FA_cout_1076;
  wire FA_cout_1077;
  wire FA_cout_1078;
  wire FA_cout_1079;
  wire FA_cout_1080;
  wire FA_cout_1081;
  wire FA_cout_1082;
  wire FA_cout_1083;
  wire FA_cout_1084;
  wire FA_cout_1085;
  wire FA_cout_1086;
  wire FA_cout_1087;
  wire FA_cout_1088;
  wire FA_cout_1089;
  wire FA_cout_1090;
  wire FA_cout_1091;
  wire FA_cout_1092;
  wire FA_cout_1093;
  wire FA_cout_1094;
  wire FA_cout_1095;
  wire FA_cout_1096;
  wire FA_cout_1097;
  wire FA_cout_1098;
  wire FA_cout_1099;
  wire FA_cout_1100;
  wire FA_cout_1101;
  wire FA_cout_1102;
  wire FA_cout_1103;
  wire FA_cout_1104;
  wire FA_cout_1105;
  wire FA_cout_1106;
  wire FA_cout_1107;
  wire FA_cout_1108;
  wire FA_cout_1109;
  wire FA_cout_1110;
  wire FA_cout_1111;
  wire FA_cout_1112;
  wire FA_cout_1113;
  wire FA_cout_1114;
  wire FA_cout_1115;
  wire FA_cout_1116;
  wire FA_cout_1117;
  wire FA_cout_1118;
  wire FA_cout_1119;
  wire FA_cout_1120;
  wire FA_cout_1121;
  wire FA_cout_1122;
  wire FA_cout_1123;
  wire FA_cout_1124;
  wire FA_cout_1125;
  wire FA_cout_1126;
  wire FA_cout_1127;
  wire FA_cout_1128;
  wire FA_cout_1129;
  wire FA_cout_1130;
  wire FA_cout_1131;
  wire FA_cout_1132;
  wire FA_cout_1133;
  wire FA_cout_1134;
  wire FA_cout_1135;
  wire FA_cout_1136;
  wire FA_cout_1137;
  wire FA_cout_1138;
  wire FA_cout_1139;
  wire FA_cout_1140;
  wire FA_cout_1141;
  wire FA_cout_1142;
  wire FA_cout_1143;
  wire FA_cout_1144;
  wire FA_cout_1145;
  wire FA_cout_1146;
  wire FA_cout_1147;
  wire FA_cout_1148;
  wire FA_cout_1149;
  wire FA_cout_1150;
  wire FA_cout_1151;
  wire FA_cout_1152;
  wire FA_cout_1153;
  wire FA_cout_1154;
  wire FA_cout_1155;
  wire FA_cout_1156;
  wire FA_cout_1157;
  wire FA_cout_1158;
  wire FA_cout_1159;
  wire FA_cout_1160;
  wire FA_cout_1161;
  wire FA_cout_1162;
  wire FA_cout_1163;
  wire FA_cout_1164;
  wire FA_cout_1165;
  wire FA_cout_1166;
  wire FA_cout_1167;
  wire FA_cout_1168;
  wire FA_cout_1169;
  wire FA_cout_1170;
  wire FA_cout_1171;
  wire FA_cout_1172;
  wire FA_cout_1173;
  wire FA_cout_1174;
  wire FA_cout_1175;
  wire FA_cout_1176;
  wire FA_cout_1177;
  wire FA_cout_1178;
  wire FA_cout_1179;
  wire FA_cout_1180;
  wire FA_cout_1181;
  wire FA_cout_1182;
  wire FA_cout_1183;
  wire FA_cout_1184;
  wire FA_cout_1185;
  wire FA_cout_1186;
  wire FA_cout_1187;
  wire FA_cout_1188;
  wire FA_cout_1189;
  wire FA_cout_1190;
  wire FA_cout_1191;
  wire FA_cout_1192;
  wire FA_cout_1193;
  wire FA_cout_1194;
  wire FA_cout_1195;
  wire FA_cout_1196;
  wire FA_cout_1197;
  wire FA_cout_1198;
  wire FA_cout_1199;
  wire FA_cout_1200;
  wire FA_cout_1201;
  wire FA_cout_1202;
  wire FA_cout_1203;
  wire FA_cout_1204;
  wire FA_cout_1205;
  wire FA_cout_1206;
  wire FA_cout_1207;
  wire FA_cout_1208;
  wire FA_cout_1209;
  wire FA_cout_1210;
  wire FA_cout_1211;
  wire FA_cout_1212;
  wire FA_cout_1213;
  wire FA_cout_1214;
  wire FA_cout_1215;
  wire FA_cout_1216;
  wire FA_cout_1217;
  wire FA_cout_1218;
  wire FA_cout_1219;
  wire FA_cout_1220;
  wire FA_cout_1221;
  wire FA_cout_1222;
  wire FA_cout_1223;
  wire FA_cout_1224;
  wire FA_cout_1225;
  wire FA_cout_1226;
  wire FA_cout_1227;
  wire FA_cout_1228;
  wire FA_cout_1229;
  wire FA_cout_1230;
  wire FA_cout_1231;
  wire FA_cout_1232;
  wire FA_cout_1233;
  wire FA_cout_1234;
  wire FA_cout_1235;
  wire FA_cout_1236;
  wire FA_cout_1237;
  wire FA_cout_1238;
  wire FA_cout_1239;
  wire FA_cout_1240;
  wire FA_cout_1241;
  wire FA_cout_1242;
  wire FA_cout_1243;
  wire FA_cout_1244;
  wire FA_cout_1245;
  wire FA_cout_1246;
  wire FA_cout_1247;
  wire FA_cout_1248;
  wire FA_cout_1249;
  wire FA_cout_1250;
  wire FA_cout_1251;
  wire FA_cout_1252;
  wire FA_cout_1253;
  wire FA_cout_1254;
  wire FA_cout_1255;
  wire FA_cout_1256;
  wire FA_cout_1257;
  wire FA_cout_1258;
  wire FA_cout_1259;
  wire FA_cout_1260;
  wire FA_cout_1261;
  wire FA_cout_1262;
  wire FA_cout_1263;
  wire FA_cout_1264;
  wire FA_cout_1265;
  wire FA_cout_1266;
  wire FA_cout_1267;
  wire FA_cout_1268;
  wire FA_cout_1269;
  wire FA_cout_1270;
  wire FA_cout_1271;
  wire FA_cout_1272;
  wire FA_cout_1273;
  wire FA_cout_1274;
  wire FA_cout_1275;
  wire FA_cout_1276;
  wire FA_cout_1277;
  wire FA_cout_1278;
  wire FA_cout_1279;
  wire FA_cout_1280;
  wire FA_cout_1281;
  wire FA_cout_1282;
  wire FA_cout_1283;
  wire FA_cout_1284;
  wire FA_cout_1285;
  wire FA_cout_1286;
  wire FA_cout_1287;
  wire FA_cout_1288;
  wire FA_cout_1289;
  wire FA_cout_1290;
  wire FA_cout_1291;
  wire FA_cout_1292;
  wire FA_cout_1293;
  wire FA_cout_1294;
  wire FA_cout_1295;
  wire FA_cout_1296;
  wire FA_cout_1297;
  wire FA_cout_1298;
  wire FA_cout_1299;
  wire FA_cout_1300;
  wire FA_cout_1301;
  wire FA_cout_1302;
  wire FA_cout_1303;
  wire FA_cout_1304;
  wire FA_cout_1305;
  wire FA_cout_1306;
  wire FA_cout_1307;
  wire FA_cout_1308;
  wire FA_cout_1309;
  wire FA_cout_1310;
  wire FA_cout_1311;
  wire FA_cout_1312;
  wire FA_cout_1313;
  wire FA_cout_1314;
  wire FA_cout_1315;
  wire FA_cout_1316;
  wire FA_cout_1317;
  wire FA_cout_1318;
  wire FA_cout_1319;
  wire FA_cout_1320;
  wire FA_cout_1321;
  wire FA_cout_1322;
  wire FA_cout_1323;
  wire FA_cout_1324;
  wire FA_cout_1325;
  wire FA_cout_1326;
  wire FA_cout_1327;
  wire FA_cout_1328;
  wire FA_cout_1329;
  wire FA_cout_1330;
  wire FA_cout_1331;
  wire FA_cout_1332;
  wire FA_cout_1333;
  wire FA_cout_1334;
  wire FA_cout_1335;
  wire FA_cout_1336;
  wire FA_cout_1337;
  wire FA_cout_1338;
  wire FA_cout_1339;
  wire FA_cout_1340;
  wire FA_cout_1341;
  wire FA_cout_1342;
  wire FA_cout_1343;
  wire FA_cout_1344;
  wire FA_cout_1345;
  wire FA_cout_1346;
  wire FA_cout_1347;
  wire FA_cout_1348;
  wire FA_cout_1349;
  wire FA_cout_1350;
  wire FA_cout_1351;
  wire FA_cout_1352;
  wire FA_cout_1353;
  wire FA_cout_1354;
  wire FA_cout_1355;
  wire FA_cout_1356;
  wire FA_cout_1357;
  wire FA_cout_1358;
  wire FA_cout_1359;
  wire FA_cout_1360;
  wire FA_cout_1361;
  wire FA_cout_1362;
  wire FA_cout_1363;
  wire FA_cout_1364;
  wire FA_cout_1365;
  wire FA_cout_1366;
  wire FA_cout_1367;
  wire FA_cout_1368;
  wire FA_cout_1369;
  wire FA_cout_1370;
  wire FA_cout_1371;
  wire FA_cout_1372;
  wire FA_cout_1373;
  wire FA_cout_1374;
  wire FA_cout_1375;
  wire FA_cout_1376;
  wire FA_cout_1377;
  wire FA_cout_1378;
  wire FA_cout_1379;
  wire FA_cout_1380;
  wire FA_cout_1381;
  wire FA_cout_1382;
  wire FA_cout_1383;
  wire FA_cout_1384;
  wire FA_cout_1385;
  wire FA_cout_1386;
  wire FA_cout_1387;
  wire FA_cout_1388;
  wire FA_cout_1389;
  wire FA_cout_1390;
  wire FA_cout_1391;
  wire FA_cout_1392;
  wire FA_cout_1393;
  wire FA_cout_1394;
  wire FA_cout_1395;
  wire FA_cout_1396;
  wire FA_cout_1397;
  wire FA_cout_1398;
  wire FA_cout_1399;
  wire FA_cout_1400;
  wire FA_cout_1401;
  wire FA_cout_1402;
  wire FA_cout_1403;
  wire FA_cout_1404;
  wire FA_cout_1405;
  wire FA_cout_1406;
  wire FA_cout_1407;
  wire FA_cout_1408;
  wire FA_cout_1409;
  wire FA_cout_1410;
  wire FA_cout_1411;
  wire FA_cout_1412;
  wire FA_cout_1413;
  wire FA_cout_1414;
  wire FA_cout_1415;
  wire FA_cout_1416;
  wire FA_cout_1417;
  wire FA_cout_1418;
  wire FA_cout_1419;
  wire FA_cout_1420;
  wire FA_cout_1421;
  wire FA_cout_1422;
  wire FA_cout_1423;
  wire FA_cout_1424;
  wire FA_cout_1425;
  wire FA_cout_1426;
  wire FA_cout_1427;
  wire FA_cout_1428;
  wire FA_cout_1429;
  wire FA_cout_1430;
  wire FA_cout_1431;
  wire FA_cout_1432;
  wire FA_cout_1433;
  wire FA_cout_1434;
  wire FA_cout_1435;
  wire FA_cout_1436;
  wire FA_cout_1437;
  wire FA_cout_1438;
  wire FA_cout_1439;
  wire FA_cout_1440;
  wire FA_cout_1441;
  wire FA_cout_1442;
  wire FA_cout_1443;
  wire FA_cout_1444;
  wire FA_cout_1445;
  wire FA_cout_1446;
  wire FA_cout_1447;
  wire FA_cout_1448;
  wire FA_cout_1449;
  wire FA_cout_1450;
  wire FA_cout_1451;
  wire FA_cout_1452;
  wire FA_cout_1453;
  wire FA_cout_1454;
  wire FA_cout_1455;
  wire FA_cout_1456;
  wire FA_cout_1457;
  wire FA_cout_1458;
  wire FA_cout_1459;
  wire FA_cout_1460;
  wire FA_cout_1461;
  wire FA_cout_1462;
  wire FA_cout_1463;
  wire FA_cout_1464;
  wire FA_cout_1465;
  wire FA_cout_1466;
  wire FA_cout_1467;
  wire FA_cout_1468;
  wire FA_cout_1469;
  wire FA_cout_1470;
  wire FA_cout_1471;
  wire FA_cout_1472;
  wire FA_cout_1473;
  wire FA_cout_1474;
  wire FA_cout_1475;
  wire FA_cout_1476;
  wire FA_cout_1477;
  wire FA_cout_1478;
  wire FA_cout_1479;
  wire FA_cout_1480;
  wire FA_cout_1481;
  wire FA_cout_1482;
  wire FA_cout_1483;
  wire FA_cout_1484;
  wire FA_cout_1485;
  wire FA_cout_1486;
  wire FA_cout_1487;
  wire FA_cout_1488;
  wire FA_cout_1489;
  wire FA_cout_1490;
  wire FA_cout_1491;
  wire FA_cout_1492;
  wire FA_cout_1493;
  wire FA_cout_1494;
  wire FA_cout_1495;
  wire FA_cout_1496;
  wire FA_cout_1497;
  wire FA_cout_1498;
  wire FA_cout_1499;
  wire FA_cout_1500;
  wire FA_cout_1501;
  wire FA_cout_1502;
  wire FA_cout_1503;
  wire FA_cout_1504;
  wire FA_cout_1505;
  wire FA_cout_1506;
  wire FA_cout_1507;
  wire FA_cout_1508;
  wire FA_cout_1509;
  wire FA_cout_1510;
  wire FA_cout_1511;
  wire FA_cout_1512;
  wire FA_cout_1513;
  wire FA_cout_1514;
  wire FA_cout_1515;
  wire FA_cout_1516;
  wire FA_cout_1517;
  wire FA_cout_1518;
  wire FA_cout_1519;
  wire FA_cout_1520;
  wire FA_cout_1521;
  wire FA_cout_1522;
  wire FA_cout_1523;
  wire FA_cout_1524;
  wire FA_cout_1525;
  wire FA_cout_1526;
  wire FA_cout_1527;
  wire FA_cout_1528;
  wire FA_cout_1529;
  wire FA_cout_1530;
  wire FA_cout_1531;
  wire FA_cout_1532;
  wire FA_cout_1533;
  wire FA_cout_1534;
  wire FA_cout_1535;
  wire FA_cout_1536;
  wire FA_cout_1537;
  wire FA_cout_1538;
  wire FA_cout_1539;
  wire FA_cout_1540;
  wire FA_cout_1541;
  wire FA_cout_1542;
  wire FA_cout_1543;
  wire FA_cout_1544;
  wire FA_cout_1545;
  wire FA_cout_1546;
  wire FA_cout_1547;
  wire FA_cout_1548;
  wire FA_cout_1549;
  wire FA_cout_1550;
  wire FA_cout_1551;
  wire FA_cout_1552;
  wire FA_cout_1553;
  wire FA_cout_1554;
  wire FA_cout_1555;
  wire FA_cout_1556;
  wire FA_cout_1557;
  wire FA_cout_1558;
  wire FA_cout_1559;
  wire FA_cout_1560;
  wire FA_cout_1561;
  wire FA_cout_1562;
  wire FA_cout_1563;
  wire FA_cout_1564;
  wire FA_cout_1565;
  wire FA_cout_1566;
  wire FA_cout_1567;
  wire FA_cout_1568;
  wire FA_cout_1569;
  wire FA_cout_1570;
  wire FA_cout_1571;
  wire FA_cout_1572;
  wire FA_cout_1573;
  wire FA_cout_1574;
  wire FA_cout_1575;
  wire FA_cout_1576;
  wire FA_cout_1577;
  wire FA_cout_1578;
  wire FA_cout_1579;
  wire FA_cout_1580;
  wire FA_cout_1581;
  wire FA_cout_1582;
  wire FA_cout_1583;
  wire FA_cout_1584;
  wire FA_cout_1585;
  wire FA_cout_1586;
  wire FA_cout_1587;
  wire FA_cout_1588;
  wire FA_cout_1589;
  wire FA_cout_1590;
  wire FA_cout_1591;
  wire FA_cout_1592;
  wire FA_cout_1593;
  wire FA_cout_1594;
  wire FA_cout_1595;
  wire FA_cout_1596;
  wire FA_cout_1597;
  wire FA_cout_1598;
  wire FA_cout_1599;
  wire FA_cout_1600;
  wire FA_cout_1601;
  wire FA_cout_1602;
  wire FA_cout_1603;
  wire FA_cout_1604;
  wire FA_cout_1605;
  wire FA_cout_1606;
  wire FA_cout_1607;
  wire FA_cout_1608;
  wire FA_cout_1609;
  wire FA_cout_1610;
  wire FA_cout_1611;
  wire FA_cout_1612;
  wire FA_cout_1613;
  wire FA_cout_1614;
  wire FA_cout_1615;
  wire FA_cout_1616;
  wire FA_cout_1617;
  wire FA_cout_1618;
  wire FA_cout_1619;
  wire FA_cout_1620;
  wire FA_cout_1621;
  wire FA_cout_1622;
  wire FA_cout_1623;
  wire FA_cout_1624;
  wire FA_cout_1625;
  wire FA_cout_1626;
  wire FA_cout_1627;
  wire FA_cout_1628;
  wire FA_cout_1629;
  wire FA_cout_1630;
  wire FA_cout_1631;
  wire FA_cout_1632;
  wire FA_cout_1633;
  wire FA_cout_1634;
  wire FA_cout_1635;
  wire FA_cout_1636;
  wire FA_cout_1637;
  wire FA_cout_1638;
  wire FA_cout_1639;
  wire FA_cout_1640;
  wire FA_cout_1641;
  wire FA_cout_1642;
  wire FA_cout_1643;
  wire FA_cout_1644;
  wire FA_cout_1645;
  wire FA_cout_1646;
  wire FA_cout_1647;
  wire FA_cout_1648;
  wire FA_cout_1649;
  wire FA_cout_1650;
  wire FA_cout_1651;
  wire FA_cout_1652;
  wire FA_cout_1653;
  wire FA_cout_1654;
  wire FA_cout_1655;
  wire FA_cout_1656;
  wire FA_cout_1657;
  wire FA_cout_1658;
  wire FA_cout_1659;
  wire FA_cout_1660;
  wire FA_cout_1661;
  wire FA_cout_1662;
  wire FA_cout_1663;
  wire FA_cout_1664;
  wire FA_cout_1665;
  wire FA_cout_1666;
  wire FA_cout_1667;
  wire FA_cout_1668;
  wire FA_cout_1669;
  wire FA_cout_1670;
  wire FA_cout_1671;
  wire FA_cout_1672;
  wire FA_cout_1673;
  wire FA_cout_1674;
  wire FA_cout_1675;
  wire FA_cout_1676;
  wire FA_cout_1677;
  wire FA_cout_1678;
  wire FA_cout_1679;
  wire FA_cout_1680;
  wire FA_cout_1681;
  wire FA_cout_1682;
  wire FA_cout_1683;
  wire FA_cout_1684;
  wire FA_cout_1685;
  wire FA_cout_1686;
  wire FA_cout_1687;
  wire FA_cout_1688;
  wire FA_cout_1689;
  wire FA_cout_1690;
  wire FA_cout_1691;
  wire FA_cout_1692;
  wire FA_cout_1693;
  wire FA_cout_1694;
  wire FA_cout_1695;
  wire FA_cout_1696;
  wire FA_cout_1697;
  wire FA_cout_1698;
  wire FA_cout_1699;
  wire FA_cout_1700;
  wire FA_cout_1701;
  wire FA_cout_1702;
  wire FA_cout_1703;
  wire FA_cout_1704;
  wire FA_cout_1705;
  wire FA_cout_1706;
  wire FA_cout_1707;
  wire FA_cout_1708;
  wire FA_cout_1709;
  wire FA_cout_1710;
  wire FA_cout_1711;
  wire FA_cout_1712;
  wire FA_cout_1713;
  wire FA_cout_1714;
  wire FA_cout_1715;
  wire FA_cout_1716;
  wire FA_cout_1717;
  wire FA_cout_1718;
  wire FA_cout_1719;
  wire FA_cout_1720;
  wire FA_cout_1721;
  wire FA_cout_1722;
  wire FA_cout_1723;
  wire FA_cout_1724;
  wire FA_cout_1725;
  wire FA_cout_1726;
  wire FA_cout_1727;
  wire FA_cout_1728;
  wire FA_cout_1729;
  wire FA_cout_1730;
  wire FA_cout_1731;
  wire FA_cout_1732;
  wire FA_cout_1733;
  wire FA_cout_1734;
  wire FA_cout_1735;
  wire FA_cout_1736;
  wire FA_cout_1737;
  wire FA_cout_1738;
  wire FA_cout_1739;
  wire FA_cout_1740;
  wire FA_cout_1741;
  wire FA_cout_1742;
  wire FA_cout_1743;
  wire FA_cout_1744;
  wire FA_cout_1745;
  wire FA_cout_1746;
  wire FA_cout_1747;
  wire FA_cout_1748;
  wire FA_cout_1749;
  wire FA_cout_1750;
  wire FA_cout_1751;
  wire FA_cout_1752;
  wire FA_cout_1753;
  wire FA_cout_1754;
  wire FA_cout_1755;
  wire FA_cout_1756;
  wire FA_cout_1757;
  wire FA_cout_1758;
  wire FA_cout_1759;
  wire FA_cout_1760;
  wire FA_cout_1761;
  wire FA_cout_1762;
  wire FA_cout_1763;
  wire FA_cout_1764;
  wire FA_cout_1765;
  wire FA_cout_1766;
  wire FA_cout_1767;
  wire FA_cout_1768;
  wire FA_cout_1769;
  wire FA_cout_1770;
  wire FA_cout_1771;
  wire FA_cout_1772;
  wire FA_cout_1773;
  wire FA_cout_1774;
  wire FA_cout_1775;
  wire FA_cout_1776;
  wire FA_cout_1777;
  wire FA_cout_1778;
  wire FA_cout_1779;
  wire FA_cout_1780;
  wire FA_cout_1781;
  wire FA_cout_1782;
  wire FA_cout_1783;
  wire FA_cout_1784;
  wire FA_cout_1785;
  wire FA_cout_1786;
  wire FA_cout_1787;
  wire FA_cout_1788;
  wire FA_cout_1789;
  wire FA_cout_1790;
  wire FA_cout_1791;
  wire FA_cout_1792;
  wire FA_cout_1793;
  wire FA_cout_1794;
  wire FA_cout_1795;
  wire FA_cout_1796;
  wire FA_cout_1797;
  wire FA_cout_1798;
  wire FA_cout_1799;
  wire FA_cout_1800;
  wire FA_cout_1801;
  wire FA_cout_1802;
  wire FA_cout_1803;
  wire FA_cout_1804;
  wire FA_cout_1805;
  wire FA_cout_1806;
  wire FA_cout_1807;
  wire FA_cout_1808;
  wire FA_cout_1809;
  wire FA_cout_1810;
  wire FA_cout_1811;
  wire FA_cout_1812;
  wire FA_cout_1813;
  wire FA_cout_1814;
  wire FA_cout_1815;
  wire FA_cout_1816;
  wire FA_cout_1817;
  wire FA_cout_1818;
  wire FA_cout_1819;
  wire FA_cout_1820;
  wire FA_cout_1821;
  wire FA_cout_1822;
  wire FA_cout_1823;
  wire FA_cout_1824;
  wire FA_cout_1825;
  wire FA_cout_1826;
  wire FA_cout_1827;
  wire FA_cout_1828;
  wire FA_cout_1829;
  wire FA_cout_1830;
  wire FA_cout_1831;
  wire FA_cout_1832;
  wire FA_cout_1833;
  wire FA_cout_1834;
  wire FA_cout_1835;
  wire FA_cout_1836;
  wire FA_cout_1837;
  wire FA_cout_1838;
  wire FA_cout_1839;
  wire FA_cout_1840;
  wire FA_cout_1841;
  wire FA_cout_1842;
  wire FA_cout_1843;
  wire FA_cout_1844;
  wire FA_cout_1845;
  wire FA_cout_1846;
  wire FA_cout_1847;
  wire FA_cout_1848;
  wire FA_cout_1849;
  wire FA_cout_1850;
  wire FA_cout_1851;
  wire FA_cout_1852;
  wire FA_cout_1853;
  wire FA_cout_1854;
  wire FA_cout_1855;
  wire FA_cout_1856;
  wire FA_cout_1857;
  wire FA_cout_1858;
  wire FA_cout_1859;
  wire FA_cout_1860;
  wire FA_cout_1861;
  wire FA_cout_1862;
  wire FA_cout_1863;
  wire FA_cout_1864;
  wire FA_cout_1865;
  wire FA_cout_1866;
  wire FA_cout_1867;
  wire FA_cout_1868;
  wire FA_cout_1869;
  wire FA_cout_1870;
  wire FA_cout_1871;
  wire FA_cout_1872;
  wire FA_cout_1873;
  wire FA_cout_1874;
  wire FA_cout_1875;
  wire FA_cout_1876;
  wire FA_cout_1877;
  wire FA_cout_1878;
  wire FA_cout_1879;
  wire FA_cout_1880;
  wire FA_cout_1881;
  wire FA_cout_1882;
  wire FA_cout_1883;
  wire FA_cout_1884;
  wire FA_cout_1885;
  wire FA_cout_1886;
  wire FA_cout_1887;
  wire FA_cout_1888;
  wire FA_cout_1889;
  wire FA_cout_1890;
  wire FA_cout_1891;
  wire FA_cout_1892;
  wire FA_cout_1893;
  wire FA_cout_1894;
  wire FA_cout_1895;
  wire FA_cout_1896;
  wire FA_cout_1897;
  wire FA_cout_1898;
  wire FA_cout_1899;
  wire FA_cout_1900;
  wire FA_cout_1901;
  wire FA_cout_1902;
  wire FA_cout_1903;
  wire FA_cout_1904;
  wire FA_cout_1905;
  wire FA_cout_1906;
  wire FA_cout_1907;
  wire FA_cout_1908;
  wire FA_cout_1909;
  wire FA_cout_1910;
  wire FA_cout_1911;
  wire FA_cout_1912;
  wire FA_cout_1913;
  wire FA_cout_1914;
  wire FA_cout_1915;
  wire FA_cout_1916;
  wire FA_cout_1917;
  wire FA_cout_1918;
  wire FA_cout_1919;
  wire FA_cout_1920;
  wire FA_cout_1921;
  wire FA_cout_1922;
  wire FA_cout_1923;
  wire FA_cout_1924;
  wire FA_cout_1925;
  wire FA_cout_1926;
  wire FA_cout_1927;
  wire FA_cout_1928;
  wire FA_cout_1929;
  wire FA_cout_1930;
  wire FA_cout_1931;
  wire FA_cout_1932;
  wire FA_cout_1933;
  wire FA_cout_1934;
  wire FA_cout_1935;
  wire FA_cout_1936;
  wire FA_cout_1937;
  wire FA_cout_1938;
  wire FA_cout_1939;
  wire FA_cout_1940;
  wire FA_cout_1941;
  wire FA_cout_1942;
  wire FA_cout_1943;
  wire FA_cout_1944;
  wire FA_cout_1945;
  wire FA_cout_1946;
  wire FA_cout_1947;
  wire FA_cout_1948;
  wire FA_cout_1949;
  wire FA_cout_1950;
  wire FA_cout_1951;
  wire FA_cout_1952;
  wire FA_cout_1953;
  wire FA_cout_1954;
  wire FA_cout_1955;
  wire FA_cout_1956;
  wire FA_cout_1957;
  wire FA_cout_1958;
  wire FA_cout_1959;
  wire FA_cout_1960;
  wire FA_cout_1961;
  wire FA_cout_1962;
  wire FA_cout_1963;
  wire FA_cout_1964;
  wire FA_cout_1965;
  wire FA_cout_1966;
  wire FA_cout_1967;
  wire FA_cout_1968;
  wire FA_cout_1969;
  wire FA_cout_1970;
  wire FA_cout_1971;
  wire FA_cout_1972;
  wire FA_cout_1973;
  wire FA_cout_1974;
  wire FA_cout_1975;
  wire FA_cout_1976;
  wire FA_cout_1977;
  wire FA_cout_1978;
  wire FA_cout_1979;
  wire FA_cout_1980;
  wire FA_cout_1981;
  wire FA_cout_1982;
  wire FA_cout_1983;
  wire FA_cout_1984;
  wire FA_cout_1985;
  wire FA_cout_1986;
  wire FA_cout_1987;
  wire FA_cout_1988;
  wire FA_cout_1989;
  wire FA_cout_1990;
  wire FA_cout_1991;
  wire FA_cout_1992;
  wire FA_cout_1993;
  wire FA_cout_1994;
  wire FA_cout_1995;
  wire FA_cout_1996;
  wire FA_cout_1997;
  wire FA_cout_1998;
  wire FA_cout_1999;
  wire FA_cout_2000;
  wire FA_cout_2001;
  wire FA_cout_2002;
  wire FA_cout_2003;
  wire FA_cout_2004;
  wire FA_cout_2005;
  wire FA_cout_2006;
  wire FA_cout_2007;
  wire FA_cout_2008;
  wire FA_cout_2009;
  wire FA_cout_2010;
  wire FA_cout_2011;
  wire FA_cout_2012;
  wire FA_cout_2013;
  wire FA_cout_2014;
  wire FA_cout_2015;
  wire FA_cout_2016;
  wire FA_cout_2017;
  wire FA_cout_2018;
  wire FA_cout_2019;
  wire FA_cout_2020;
  wire FA_cout_2021;
  wire FA_cout_2022;
  wire FA_cout_2023;
  wire FA_cout_2024;
  wire FA_cout_2025;
  wire FA_cout_2026;
  wire FA_cout_2027;
  wire FA_cout_2028;
  wire FA_cout_2029;
  wire FA_cout_2030;
  wire FA_cout_2031;
  wire FA_cout_2032;
  wire FA_cout_2033;
  wire FA_cout_2034;
  wire FA_cout_2035;
  wire FA_cout_2036;
  wire FA_cout_2037;
  wire FA_cout_2038;
  wire FA_cout_2039;
  wire FA_cout_2040;
  wire FA_cout_2041;
  wire FA_cout_2042;
  wire FA_cout_2043;
  wire FA_cout_2044;
  wire FA_cout_2045;
  wire FA_cout_2046;
  wire FA_cout_2047;
  wire FA_cout_2048;
  wire FA_cout_2049;
  wire FA_cout_2050;
  wire FA_cout_2051;
  wire FA_cout_2052;
  wire FA_cout_2053;
  wire FA_cout_2054;
  wire FA_cout_2055;
  wire FA_cout_2056;
  wire FA_cout_2057;
  wire FA_cout_2058;
  wire FA_cout_2059;
  wire FA_cout_2060;
  wire FA_cout_2061;
  wire FA_cout_2062;
  wire FA_cout_2063;
  wire FA_cout_2064;
  wire FA_cout_2065;
  wire FA_cout_2066;
  wire FA_cout_2067;
  wire FA_cout_2068;
  wire FA_cout_2069;
  wire FA_cout_2070;
  wire FA_cout_2071;
  wire FA_cout_2072;
  wire FA_cout_2073;
  wire FA_cout_2074;
  wire FA_cout_2075;
  wire FA_cout_2076;
  wire FA_cout_2077;
  wire FA_cout_2078;
  wire FA_cout_2079;
  wire FA_cout_2080;
  wire FA_cout_2081;
  wire FA_cout_2082;
  wire FA_cout_2083;
  wire FA_cout_2084;
  wire FA_cout_2085;
  wire FA_cout_2086;
  wire FA_cout_2087;
  wire FA_cout_2088;
  wire FA_cout_2089;
  wire FA_cout_2090;
  wire FA_cout_2091;
  wire FA_cout_2092;
  wire FA_cout_2093;
  wire FA_cout_2094;
  wire FA_cout_2095;
  wire FA_cout_2096;
  wire FA_cout_2097;
  wire FA_cout_2098;
  wire FA_cout_2099;
  wire FA_cout_2100;
  wire FA_cout_2101;
  wire FA_cout_2102;
  wire FA_cout_2103;
  wire FA_cout_2104;
  wire FA_cout_2105;
  wire FA_cout_2106;
  wire FA_cout_2107;
  wire FA_cout_2108;
  wire FA_cout_2109;
  wire FA_cout_2110;
  wire FA_cout_2111;
  wire FA_cout_2112;
  wire FA_cout_2113;
  wire FA_cout_2114;
  wire FA_cout_2115;
  wire FA_cout_2116;
  wire FA_cout_2117;
  wire FA_cout_2118;
  wire FA_cout_2119;
  wire FA_cout_2120;
  wire FA_cout_2121;
  wire FA_cout_2122;
  wire FA_cout_2123;
  wire FA_cout_2124;
  wire FA_cout_2125;
  wire FA_cout_2126;
  wire FA_cout_2127;
  wire FA_cout_2128;
  wire FA_cout_2129;
  wire FA_cout_2130;
  wire FA_cout_2131;
  wire FA_cout_2132;
  wire FA_cout_2133;
  wire FA_cout_2134;
  wire FA_cout_2135;
  wire FA_cout_2136;
  wire FA_cout_2137;
  wire FA_cout_2138;
  wire FA_cout_2139;
  wire FA_cout_2140;
  wire FA_cout_2141;
  wire FA_cout_2142;
  wire FA_cout_2143;
  wire FA_cout_2144;
  wire FA_cout_2145;
  wire FA_cout_2146;
  wire FA_cout_2147;
  wire FA_cout_2148;
  wire FA_cout_2149;
  wire FA_cout_2150;
  wire FA_cout_2151;
  wire FA_cout_2152;
  wire FA_cout_2153;
  wire FA_cout_2154;
  wire FA_cout_2155;
  wire FA_cout_2156;
  wire FA_cout_2157;
  wire FA_cout_2158;
  wire FA_cout_2159;
  wire FA_cout_2160;
  wire FA_cout_2161;
  wire FA_cout_2162;
  wire FA_cout_2163;
  wire FA_cout_2164;
  wire FA_cout_2165;
  wire FA_cout_2166;
  wire FA_cout_2167;
  wire FA_cout_2168;
  wire FA_cout_2169;
  wire FA_cout_2170;
  wire FA_cout_2171;
  wire FA_cout_2172;
  wire FA_cout_2173;
  wire FA_cout_2174;
  wire FA_cout_2175;
  wire FA_cout_2176;
  wire FA_cout_2177;
  wire FA_cout_2178;
  wire FA_cout_2179;
  wire FA_cout_2180;
  wire FA_cout_2181;
  wire FA_cout_2182;
  wire FA_cout_2183;
  wire FA_cout_2184;
  wire FA_cout_2185;
  wire FA_cout_2186;
  wire FA_cout_2187;
  wire FA_cout_2188;
  wire FA_cout_2189;
  wire FA_cout_2190;
  wire FA_cout_2191;
  wire FA_cout_2192;
  wire FA_cout_2193;
  wire FA_cout_2194;
  wire FA_cout_2195;
  wire FA_cout_2196;
  wire FA_cout_2197;
  wire FA_cout_2198;
  wire FA_cout_2199;
  wire FA_cout_2200;
  wire FA_cout_2201;
  wire FA_cout_2202;
  wire FA_cout_2203;
  wire FA_cout_2204;
  wire FA_cout_2205;
  wire FA_cout_2206;
  wire FA_cout_2207;
  wire FA_cout_2208;
  wire FA_cout_2209;
  wire FA_cout_2210;
  wire FA_cout_2211;
  wire FA_cout_2212;
  wire FA_cout_2213;
  wire FA_cout_2214;
  wire FA_cout_2215;
  wire FA_cout_2216;
  wire FA_cout_2217;
  wire FA_cout_2218;
  wire FA_cout_2219;
  wire FA_cout_2220;
  wire FA_cout_2221;
  wire FA_cout_2222;
  wire FA_cout_2223;
  wire FA_cout_2224;
  wire FA_cout_2225;
  wire FA_cout_2226;
  wire FA_cout_2227;
  wire FA_cout_2228;
  wire FA_cout_2229;
  wire FA_cout_2230;
  wire FA_cout_2231;
  wire FA_cout_2232;
  wire FA_cout_2233;
  wire FA_cout_2234;
  wire FA_cout_2235;
  wire FA_cout_2236;
  wire FA_cout_2237;
  wire FA_cout_2238;
  wire FA_cout_2239;
  wire FA_cout_2240;
  wire FA_cout_2241;
  wire FA_cout_2242;
  wire FA_cout_2243;
  wire FA_cout_2244;
  wire FA_cout_2245;
  wire FA_cout_2246;
  wire FA_cout_2247;
  wire FA_cout_2248;
  wire FA_cout_2249;
  wire FA_cout_2250;
  wire FA_cout_2251;
  wire FA_cout_2252;
  wire FA_cout_2253;
  wire FA_cout_2254;
  wire FA_cout_2255;
  wire FA_cout_2256;
  wire FA_cout_2257;
  wire FA_cout_2258;
  wire FA_cout_2259;
  wire FA_cout_2260;
  wire FA_cout_2261;
  wire FA_cout_2262;
  wire FA_cout_2263;
  wire FA_cout_2264;
  wire FA_cout_2265;
  wire FA_cout_2266;
  wire FA_cout_2267;
  wire FA_cout_2268;
  wire FA_cout_2269;
  wire FA_cout_2270;
  wire FA_cout_2271;
  wire FA_cout_2272;
  wire FA_cout_2273;
  wire FA_cout_2274;
  wire FA_cout_2275;
  wire FA_cout_2276;
  wire FA_cout_2277;
  wire FA_cout_2278;
  wire FA_cout_2279;
  wire FA_cout_2280;
  wire FA_cout_2281;
  wire FA_cout_2282;
  wire FA_cout_2283;
  wire FA_cout_2284;
  wire FA_cout_2285;
  wire FA_cout_2286;
  wire FA_cout_2287;
  wire FA_cout_2288;
  wire FA_cout_2289;
  wire FA_cout_2290;
  wire FA_cout_2291;
  wire FA_cout_2292;
  wire FA_cout_2293;
  wire FA_cout_2294;
  wire FA_cout_2295;
  wire FA_cout_2296;
  wire FA_cout_2297;
  wire FA_cout_2298;
  wire FA_cout_2299;
  wire FA_cout_2300;
  wire FA_cout_2301;
  wire FA_cout_2302;
  wire FA_cout_2303;
  wire FA_cout_2304;
  wire FA_cout_2305;
  wire FA_cout_2306;
  wire FA_cout_2307;
  wire FA_cout_2308;
  wire FA_cout_2309;
  wire FA_cout_2310;
  wire FA_cout_2311;
  wire FA_cout_2312;
  wire FA_cout_2313;
  wire FA_cout_2314;
  wire FA_cout_2315;
  wire FA_cout_2316;
  wire FA_cout_2317;
  wire FA_cout_2318;
  wire FA_cout_2319;
  wire FA_cout_2320;
  wire FA_cout_2321;
  wire FA_cout_2322;
  wire FA_cout_2323;
  wire FA_cout_2324;
  wire FA_cout_2325;
  wire FA_cout_2326;
  wire FA_cout_2327;
  wire FA_cout_2328;
  wire FA_cout_2329;
  wire FA_cout_2330;
  wire FA_cout_2331;
  wire FA_cout_2332;
  wire FA_cout_2333;
  wire FA_cout_2334;
  wire FA_cout_2335;
  wire FA_cout_2336;
  wire FA_cout_2337;
  wire FA_cout_2338;
  wire FA_cout_2339;
  wire FA_cout_2340;
  wire FA_cout_2341;
  wire FA_cout_2342;
  wire FA_cout_2343;
  wire FA_cout_2344;
  wire FA_cout_2345;
  wire FA_cout_2346;
  wire FA_cout_2347;
  wire FA_cout_2348;
  wire FA_cout_2349;
  wire FA_cout_2350;
  wire FA_cout_2351;
  wire FA_cout_2352;
  wire FA_cout_2353;
  wire FA_cout_2354;
  wire FA_cout_2355;
  wire FA_cout_2356;
  wire FA_cout_2357;
  wire FA_cout_2358;
  wire FA_cout_2359;
  wire FA_cout_2360;
  wire FA_cout_2361;
  wire FA_cout_2362;
  wire FA_cout_2363;
  wire FA_cout_2364;
  wire FA_cout_2365;
  wire FA_cout_2366;
  wire FA_cout_2367;
  wire FA_cout_2368;
  wire FA_cout_2369;
  wire FA_cout_2370;
  wire FA_cout_2371;
  wire FA_cout_2372;
  wire FA_cout_2373;
  wire FA_cout_2374;
  wire FA_cout_2375;
  wire FA_cout_2376;
  wire FA_cout_2377;
  wire FA_cout_2378;
  wire FA_cout_2379;
  wire FA_cout_2380;
  wire FA_cout_2381;
  wire FA_cout_2382;
  wire FA_cout_2383;
  wire FA_cout_2384;
  wire FA_cout_2385;
  wire FA_cout_2386;
  wire FA_cout_2387;
  wire FA_cout_2388;
  wire FA_cout_2389;
  wire FA_cout_2390;
  wire FA_cout_2391;
  wire FA_cout_2392;
  wire FA_cout_2393;
  wire FA_cout_2394;
  wire FA_cout_2395;
  wire FA_cout_2396;
  wire FA_cout_2397;
  wire FA_cout_2398;
  wire FA_cout_2399;
  wire FA_cout_2400;
  wire FA_cout_2401;
  wire FA_cout_2402;
  wire FA_cout_2403;
  wire FA_cout_2404;
  wire FA_cout_2405;
  wire FA_cout_2406;
  wire FA_cout_2407;
  wire FA_cout_2408;
  wire FA_cout_2409;
  wire FA_cout_2410;
  wire FA_cout_2411;
  wire FA_cout_2412;
  wire FA_cout_2413;
  wire FA_cout_2414;
  wire FA_cout_2415;
  wire FA_cout_2416;
  wire FA_cout_2417;
  wire FA_cout_2418;
  wire FA_cout_2419;
  wire FA_cout_2420;
  wire FA_cout_2421;
  wire FA_cout_2422;
  wire FA_cout_2423;
  wire FA_cout_2424;
  wire FA_cout_2425;
  wire FA_cout_2426;
  wire FA_cout_2427;
  wire FA_cout_2428;
  wire FA_cout_2429;
  wire FA_cout_2430;
  wire FA_cout_2431;
  wire FA_cout_2432;
  wire FA_cout_2433;
  wire FA_cout_2434;
  wire FA_cout_2435;
  wire FA_cout_2436;
  wire FA_cout_2437;
  wire FA_cout_2438;
  wire FA_cout_2439;
  wire FA_cout_2440;
  wire FA_cout_2441;
  wire FA_cout_2442;
  wire FA_cout_2443;
  wire FA_cout_2444;
  wire FA_cout_2445;
  wire FA_cout_2446;
  wire FA_cout_2447;
  wire FA_cout_2448;
  wire FA_cout_2449;
  wire FA_cout_2450;
  wire FA_cout_2451;
  wire FA_cout_2452;
  wire FA_cout_2453;
  wire FA_cout_2454;
  wire FA_cout_2455;
  wire FA_cout_2456;
  wire FA_cout_2457;
  wire FA_cout_2458;
  wire FA_cout_2459;
  wire FA_cout_2460;
  wire FA_cout_2461;
  wire FA_cout_2462;
  wire FA_cout_2463;
  wire FA_cout_2464;
  wire FA_cout_2465;
  wire FA_cout_2466;
  wire FA_cout_2467;
  wire FA_cout_2468;
  wire FA_cout_2469;
  wire FA_cout_2470;
  wire FA_cout_2471;
  wire FA_cout_2472;
  wire FA_cout_2473;
  wire FA_cout_2474;
  wire FA_cout_2475;
  wire FA_cout_2476;
  wire FA_cout_2477;
  wire FA_cout_2478;
  wire FA_cout_2479;
  wire FA_cout_2480;
  wire FA_cout_2481;
  wire FA_cout_2482;
  wire FA_cout_2483;
  wire FA_cout_2484;
  wire FA_cout_2485;
  wire FA_cout_2486;
  wire FA_cout_2487;
  wire FA_cout_2488;
  wire FA_cout_2489;
  wire FA_cout_2490;
  wire FA_cout_2491;
  wire FA_cout_2492;
  wire FA_cout_2493;
  wire FA_cout_2494;
  wire FA_cout_2495;
  wire FA_cout_2496;
  wire FA_cout_2497;
  wire FA_cout_2498;
  wire FA_cout_2499;
  wire FA_cout_2500;
  wire FA_cout_2501;
  wire FA_cout_2502;
  wire FA_cout_2503;
  wire FA_cout_2504;
  wire FA_cout_2505;
  wire FA_cout_2506;
  wire FA_cout_2507;
  wire FA_cout_2508;
  wire FA_cout_2509;
  wire FA_cout_2510;
  wire FA_cout_2511;
  wire FA_cout_2512;
  wire FA_cout_2513;
  wire FA_cout_2514;
  wire FA_cout_2515;
  wire FA_cout_2516;
  wire FA_cout_2517;
  wire FA_cout_2518;
  wire FA_cout_2519;
  wire FA_cout_2520;
  wire FA_cout_2521;
  wire FA_cout_2522;
  wire FA_cout_2523;
  wire FA_cout_2524;
  wire FA_cout_2525;
  wire FA_cout_2526;
  wire FA_cout_2527;
  wire FA_cout_2528;
  wire FA_cout_2529;
  wire FA_cout_2530;
  wire FA_cout_2531;
  wire FA_cout_2532;
  wire FA_cout_2533;
  wire FA_cout_2534;
  wire FA_cout_2535;
  wire FA_cout_2536;
  wire FA_cout_2537;
  wire FA_cout_2538;
  wire FA_cout_2539;
  wire FA_cout_2540;
  wire FA_cout_2541;
  wire FA_cout_2542;
  wire FA_cout_2543;
  wire FA_cout_2544;
  wire FA_cout_2545;
  wire FA_cout_2546;
  wire FA_cout_2547;
  wire FA_cout_2548;
  wire FA_cout_2549;
  wire FA_cout_2550;
  wire FA_cout_2551;
  wire FA_cout_2552;
  wire FA_cout_2553;
  wire FA_cout_2554;
  wire FA_cout_2555;
  wire FA_cout_2556;
  wire FA_cout_2557;
  wire FA_cout_2558;
  wire FA_cout_2559;
  wire FA_cout_2560;
  wire FA_cout_2561;
  wire FA_cout_2562;
  wire FA_cout_2563;
  wire FA_cout_2564;
  wire FA_cout_2565;
  wire FA_cout_2566;
  wire FA_cout_2567;
  wire FA_cout_2568;
  wire FA_cout_2569;
  wire FA_cout_2570;
  wire FA_cout_2571;
  wire FA_cout_2572;
  wire FA_cout_2573;
  wire FA_cout_2574;
  wire FA_cout_2575;
  wire FA_cout_2576;
  wire FA_cout_2577;
  wire FA_cout_2578;
  wire FA_cout_2579;
  wire FA_cout_2580;
  wire FA_cout_2581;
  wire FA_cout_2582;
  wire FA_cout_2583;
  wire FA_cout_2584;
  wire FA_cout_2585;
  wire FA_cout_2586;
  wire FA_cout_2587;
  wire FA_cout_2588;
  wire FA_cout_2589;
  wire FA_cout_2590;
  wire FA_cout_2591;
  wire FA_cout_2592;
  wire FA_cout_2593;
  wire FA_cout_2594;
  wire FA_cout_2595;
  wire FA_cout_2596;
  wire FA_cout_2597;
  wire FA_cout_2598;
  wire FA_cout_2599;
  wire FA_cout_2600;
  wire FA_cout_2601;
  wire FA_cout_2602;
  wire FA_cout_2603;
  wire FA_cout_2604;
  wire FA_cout_2605;
  wire FA_cout_2606;
  wire FA_cout_2607;
  wire FA_cout_2608;
  wire FA_cout_2609;
  wire FA_cout_2610;
  wire FA_cout_2611;
  wire FA_cout_2612;
  wire FA_cout_2613;
  wire FA_cout_2614;
  wire FA_cout_2615;
  wire FA_cout_2616;
  wire FA_cout_2617;
  wire FA_cout_2618;
  wire FA_cout_2619;
  wire FA_cout_2620;
  wire FA_cout_2621;
  wire FA_cout_2622;
  wire FA_cout_2623;
  wire FA_cout_2624;
  wire FA_cout_2625;
  wire FA_cout_2626;
  wire FA_cout_2627;
  wire FA_cout_2628;
  wire FA_cout_2629;
  wire FA_cout_2630;
  wire FA_cout_2631;
  wire FA_cout_2632;
  wire FA_cout_2633;
  wire FA_cout_2634;
  wire FA_cout_2635;
  wire FA_cout_2636;
  wire FA_cout_2637;
  wire FA_cout_2638;
  wire FA_cout_2639;
  wire FA_cout_2640;
  wire FA_cout_2641;
  wire FA_cout_2642;
  wire FA_cout_2643;
  wire FA_cout_2644;
  wire FA_cout_2645;
  wire FA_cout_2646;
  wire FA_cout_2647;
  wire FA_cout_2648;
  wire FA_cout_2649;
  wire FA_cout_2650;
  wire FA_cout_2651;
  wire FA_cout_2652;
  wire FA_cout_2653;
  wire FA_cout_2654;
  wire FA_cout_2655;
  wire FA_cout_2656;
  wire FA_cout_2657;
  wire FA_cout_2658;
  wire FA_cout_2659;
  wire FA_cout_2660;
  wire FA_cout_2661;
  wire FA_cout_2662;
  wire FA_cout_2663;
  wire FA_cout_2664;
  wire FA_cout_2665;
  wire FA_cout_2666;
  wire FA_cout_2667;
  wire FA_cout_2668;
  wire FA_cout_2669;
  wire FA_cout_2670;
  wire FA_cout_2671;
  wire FA_cout_2672;
  wire FA_cout_2673;
  wire FA_cout_2674;
  wire FA_cout_2675;
  wire FA_cout_2676;
  wire FA_cout_2677;
  wire FA_cout_2678;
  wire FA_cout_2679;
  wire FA_cout_2680;
  wire FA_cout_2681;
  wire FA_cout_2682;
  wire FA_cout_2683;
  wire FA_cout_2684;
  wire FA_cout_2685;
  wire FA_cout_2686;
  wire FA_cout_2687;
  wire FA_cout_2688;
  wire FA_cout_2689;
  wire FA_cout_2690;
  wire FA_cout_2691;
  wire FA_cout_2692;
  wire FA_cout_2693;
  wire FA_cout_2694;
  wire FA_cout_2695;
  wire FA_cout_2696;
  wire FA_cout_2697;
  wire FA_cout_2698;
  wire FA_cout_2699;
  wire FA_cout_2700;
  wire FA_cout_2701;
  wire FA_cout_2702;
  wire FA_cout_2703;
  wire FA_cout_2704;
  wire FA_cout_2705;
  wire FA_cout_2706;
  wire FA_cout_2707;
  wire FA_cout_2708;
  wire FA_cout_2709;
  wire FA_cout_2710;
  wire FA_cout_2711;
  wire FA_cout_2712;
  wire FA_cout_2713;
  wire FA_cout_2714;
  wire FA_cout_2715;
  wire FA_cout_2716;
  wire FA_cout_2717;
  wire FA_cout_2718;
  wire FA_cout_2719;
  wire FA_cout_2720;
  wire FA_cout_2721;
  wire FA_cout_2722;
  wire FA_cout_2723;
  wire FA_cout_2724;
  wire FA_cout_2725;
  wire FA_cout_2726;
  wire FA_cout_2727;
  wire FA_cout_2728;
  wire FA_cout_2729;
  wire FA_cout_2730;
  wire FA_cout_2731;
  wire FA_cout_2732;
  wire FA_cout_2733;
  wire FA_cout_2734;
  wire FA_cout_2735;
  wire FA_cout_2736;
  wire FA_cout_2737;
  wire FA_cout_2738;
  wire FA_cout_2739;
  wire FA_cout_2740;
  wire FA_cout_2741;
  wire FA_cout_2742;
  wire FA_cout_2743;
  wire FA_cout_2744;
  wire FA_cout_2745;
  wire FA_cout_2746;
  wire FA_cout_2747;
  wire FA_cout_2748;
  wire FA_cout_2749;
  wire FA_cout_2750;
  wire FA_cout_2751;
  wire FA_cout_2752;
  wire FA_cout_2753;
  wire FA_cout_2754;
  wire FA_cout_2755;
  wire FA_cout_2756;
  wire FA_cout_2757;
  wire FA_cout_2758;
  wire FA_cout_2759;
  wire FA_cout_2760;
  wire FA_cout_2761;
  wire FA_cout_2762;
  wire FA_cout_2763;
  wire FA_cout_2764;
  wire FA_cout_2765;
  wire FA_cout_2766;
  wire FA_cout_2767;
  wire FA_cout_2768;
  wire FA_cout_2769;
  wire FA_cout_2770;
  wire FA_cout_2771;
  wire FA_cout_2772;
  wire FA_cout_2773;
  wire FA_cout_2774;
  wire FA_cout_2775;
  wire FA_cout_2776;
  wire FA_cout_2777;
  wire FA_cout_2778;
  wire FA_cout_2779;
  wire FA_cout_2780;
  wire FA_cout_2781;
  wire FA_cout_2782;
  wire FA_cout_2783;
  wire FA_cout_2784;
  wire FA_cout_2785;
  wire FA_cout_2786;
  wire FA_cout_2787;
  wire FA_cout_2788;
  wire FA_cout_2789;
  wire FA_cout_2790;
  wire FA_cout_2791;
  wire FA_cout_2792;
  wire FA_cout_2793;
  wire FA_cout_2794;
  wire FA_cout_2795;
  wire FA_cout_2796;
  wire FA_cout_2797;
  wire FA_cout_2798;
  wire FA_cout_2799;
  wire FA_cout_2800;
  wire FA_cout_2801;
  wire FA_cout_2802;
  wire FA_cout_2803;
  wire FA_cout_2804;
  wire FA_cout_2805;
  wire FA_cout_2806;
  wire FA_cout_2807;
  wire FA_cout_2808;
  wire FA_cout_2809;
  wire FA_cout_2810;
  wire FA_cout_2811;
  wire FA_cout_2812;
  wire FA_cout_2813;
  wire FA_cout_2814;
  wire FA_cout_2815;
  wire FA_cout_2816;
  wire FA_cout_2817;
  wire FA_cout_2818;
  wire FA_cout_2819;
  wire FA_cout_2820;
  wire FA_cout_2821;
  wire FA_cout_2822;
  wire FA_cout_2823;
  wire FA_cout_2824;
  wire FA_cout_2825;
  wire FA_cout_2826;
  wire FA_cout_2827;
  wire FA_cout_2828;
  wire FA_cout_2829;
  wire FA_cout_2830;
  wire FA_cout_2831;
  wire FA_cout_2832;
  wire FA_cout_2833;
  wire FA_cout_2834;
  wire FA_cout_2835;
  wire FA_cout_2836;
  wire FA_cout_2837;
  wire FA_cout_2838;
  wire FA_cout_2839;
  wire FA_cout_2840;
  wire FA_cout_2841;
  wire FA_cout_2842;
  wire FA_cout_2843;
  wire FA_cout_2844;
  wire FA_cout_2845;
  wire FA_cout_2846;
  wire FA_cout_2847;
  wire FA_cout_2848;
  wire FA_cout_2849;
  wire FA_cout_2850;
  wire FA_cout_2851;
  wire FA_cout_2852;
  wire FA_cout_2853;
  wire FA_cout_2854;
  wire FA_cout_2855;
  wire FA_cout_2856;
  wire FA_cout_2857;
  wire FA_cout_2858;
  wire FA_cout_2859;
  wire FA_cout_2860;
  wire FA_cout_2861;
  wire FA_cout_2862;
  wire FA_cout_2863;
  wire FA_cout_2864;
  wire FA_cout_2865;
  wire FA_cout_2866;
  wire FA_cout_2867;
  wire FA_cout_2868;
  wire FA_cout_2869;
  wire FA_cout_2870;
  wire FA_cout_2871;
  wire FA_cout_2872;
  wire FA_cout_2873;
  wire FA_cout_2874;
  wire FA_cout_2875;
  wire FA_cout_2876;
  wire FA_cout_2877;
  wire FA_cout_2878;
  wire FA_cout_2879;
  wire FA_cout_2880;
  wire FA_cout_2881;
  wire FA_cout_2882;
  wire FA_cout_2883;
  wire FA_cout_2884;
  wire FA_cout_2885;
  wire FA_cout_2886;
  wire FA_cout_2887;
  wire FA_cout_2888;
  wire FA_cout_2889;
  wire FA_cout_2890;
  wire FA_cout_2891;
  wire FA_cout_2892;
  wire FA_cout_2893;
  wire FA_cout_2894;
  wire FA_cout_2895;
  wire FA_cout_2896;
  wire FA_cout_2897;
  wire FA_cout_2898;
  wire FA_cout_2899;
  wire FA_cout_2900;
  wire FA_cout_2901;
  wire FA_cout_2902;
  wire FA_cout_2903;
  wire FA_cout_2904;
  wire FA_cout_2905;
  wire FA_cout_2906;
  wire FA_cout_2907;
  wire FA_cout_2908;
  wire FA_cout_2909;
  wire FA_cout_2910;
  wire FA_cout_2911;
  wire FA_cout_2912;
  wire FA_cout_2913;
  wire FA_cout_2914;
  wire FA_cout_2915;
  wire FA_cout_2916;
  wire FA_cout_2917;
  wire FA_cout_2918;
  wire FA_cout_2919;
  wire FA_cout_2920;
  wire FA_cout_2921;
  wire FA_cout_2922;
  wire FA_cout_2923;
  wire FA_cout_2924;
  wire FA_cout_2925;
  wire FA_cout_2926;
  wire FA_cout_2927;
  wire FA_cout_2928;
  wire FA_cout_2929;
  wire FA_cout_2930;
  wire FA_cout_2931;
  wire FA_cout_2932;
  wire FA_cout_2933;
  wire FA_cout_2934;
  wire FA_cout_2935;
  wire FA_cout_2936;
  wire FA_cout_2937;
  wire FA_cout_2938;
  wire FA_cout_2939;
  wire FA_cout_2940;
  wire FA_cout_2941;
  wire FA_cout_2942;
  wire FA_cout_2943;
  wire FA_cout_2944;
  wire FA_cout_2945;
  wire FA_cout_2946;
  wire FA_cout_2947;
  wire FA_cout_2948;
  wire FA_cout_2949;
  wire FA_cout_2950;
  wire FA_cout_2951;
  wire FA_cout_2952;
  wire FA_cout_2953;
  wire FA_cout_2954;
  wire FA_cout_2955;
  wire FA_cout_2956;
  wire FA_cout_2957;
  wire FA_cout_2958;
  wire FA_cout_2959;
  wire FA_cout_2960;
  wire FA_cout_2961;
  wire FA_cout_2962;
  wire FA_cout_2963;
  wire FA_cout_2964;
  wire FA_cout_2965;
  wire FA_cout_2966;
  wire FA_cout_2967;
  wire FA_cout_2968;
  wire FA_cout_2969;
  wire FA_cout_2970;
  wire FA_cout_2971;
  wire FA_cout_2972;
  wire FA_cout_2973;
  wire FA_cout_2974;
  wire FA_cout_2975;
  wire FA_cout_2976;
  wire FA_cout_2977;
  wire FA_cout_2978;
  wire FA_cout_2979;
  wire FA_cout_2980;
  wire FA_cout_2981;
  wire FA_cout_2982;
  wire FA_cout_2983;
  wire FA_cout_2984;
  wire FA_cout_2985;
  wire FA_cout_2986;
  wire FA_cout_2987;
  wire FA_cout_2988;
  wire FA_cout_2989;
  wire FA_cout_2990;
  wire FA_cout_2991;
  wire FA_cout_2992;
  wire FA_cout_2993;
  wire FA_cout_2994;
  wire FA_cout_2995;
  wire FA_cout_2996;
  wire FA_cout_2997;
  wire FA_cout_2998;
  wire FA_cout_2999;
  wire FA_cout_3000;
  wire FA_cout_3001;
  wire FA_cout_3002;
  wire FA_cout_3003;
  wire FA_cout_3004;
  wire FA_cout_3005;
  wire FA_cout_3006;
  wire FA_cout_3007;
  wire FA_cout_3008;
  wire FA_cout_3009;
  wire FA_cout_3010;
  wire FA_cout_3011;
  wire FA_cout_3012;
  wire FA_cout_3013;
  wire FA_cout_3014;
  wire FA_cout_3015;
  wire FA_cout_3016;
  wire FA_cout_3017;
  wire FA_cout_3018;
  wire FA_cout_3019;
  wire FA_cout_3020;
  wire FA_cout_3021;
  wire FA_cout_3022;
  wire FA_cout_3023;
  wire FA_cout_3024;
  wire FA_cout_3025;
  wire FA_cout_3026;
  wire FA_cout_3027;
  wire FA_cout_3028;
  wire FA_cout_3029;
  wire FA_cout_3030;
  wire FA_cout_3031;
  wire FA_cout_3032;
  wire FA_cout_3033;
  wire FA_cout_3034;
  wire FA_cout_3035;
  wire FA_cout_3036;
  wire FA_cout_3037;
  wire FA_cout_3038;
  wire FA_cout_3039;
  wire FA_cout_3040;
  wire FA_cout_3041;
  wire FA_cout_3042;
  wire FA_cout_3043;
  wire FA_cout_3044;
  wire FA_cout_3045;
  wire FA_cout_3046;
  wire FA_cout_3047;
  wire FA_cout_3048;
  wire FA_cout_3049;
  wire FA_cout_3050;
  wire FA_cout_3051;
  wire FA_cout_3052;
  wire FA_cout_3053;
  wire FA_cout_3054;
  wire FA_cout_3055;
  wire FA_cout_3056;
  wire FA_cout_3057;
  wire FA_cout_3058;
  wire FA_cout_3059;
  wire FA_cout_3060;
  wire FA_cout_3061;
  wire FA_cout_3062;
  wire FA_cout_3063;
  wire FA_cout_3064;
  wire FA_cout_3065;
  wire FA_cout_3066;
  wire FA_cout_3067;
  wire FA_cout_3068;
  wire FA_cout_3069;
  wire FA_cout_3070;
  wire FA_cout_3071;
  wire FA_cout_3072;
  wire FA_cout_3073;
  wire FA_cout_3074;
  wire FA_cout_3075;
  wire FA_cout_3076;
  wire FA_cout_3077;
  wire FA_cout_3078;
  wire FA_cout_3079;
  wire FA_cout_3080;
  wire FA_cout_3081;
  wire FA_cout_3082;
  wire FA_cout_3083;
  wire FA_cout_3084;
  wire FA_cout_3085;
  wire FA_cout_3086;
  wire FA_cout_3087;
  wire FA_cout_3088;
  wire FA_cout_3089;
  wire FA_cout_3090;
  wire FA_cout_3091;
  wire FA_cout_3092;
  wire FA_cout_3093;
  wire FA_cout_3094;
  wire FA_cout_3095;
  wire FA_cout_3096;
  wire FA_cout_3097;
  wire FA_cout_3098;
  wire FA_cout_3099;
  wire FA_cout_3100;
  wire FA_cout_3101;
  wire FA_cout_3102;
  wire FA_cout_3103;
  wire FA_cout_3104;
  wire FA_cout_3105;
  wire FA_cout_3106;
  wire FA_cout_3107;
  wire FA_cout_3108;
  wire FA_cout_3109;
  wire FA_cout_3110;
  wire FA_cout_3111;
  wire FA_cout_3112;
  wire FA_cout_3113;
  wire FA_cout_3114;
  wire FA_cout_3115;
  wire FA_cout_3116;
  wire FA_cout_3117;
  wire FA_cout_3118;
  wire FA_cout_3119;
  wire FA_cout_3120;
  wire FA_cout_3121;
  wire FA_cout_3122;
  wire FA_cout_3123;
  wire FA_cout_3124;
  wire FA_cout_3125;
  wire FA_cout_3126;
  wire FA_cout_3127;
  wire FA_cout_3128;
  wire FA_cout_3129;
  wire FA_cout_3130;
  wire FA_cout_3131;
  wire FA_cout_3132;
  wire FA_cout_3133;
  wire FA_cout_3134;
  wire FA_cout_3135;
  wire FA_cout_3136;
  wire FA_cout_3137;
  wire FA_cout_3138;
  wire FA_cout_3139;
  wire FA_cout_3140;
  wire FA_cout_3141;
  wire FA_cout_3142;
  wire FA_cout_3143;
  wire FA_cout_3144;
  wire FA_cout_3145;
  wire FA_cout_3146;
  wire FA_cout_3147;
  wire FA_cout_3148;
  wire FA_cout_3149;
  wire FA_cout_3150;
  wire FA_cout_3151;
  wire FA_cout_3152;
  wire FA_cout_3153;
  wire FA_cout_3154;
  wire FA_cout_3155;
  wire FA_cout_3156;
  wire FA_cout_3157;
  wire FA_cout_3158;
  wire FA_cout_3159;
  wire FA_cout_3160;
  wire FA_cout_3161;
  wire FA_cout_3162;
  wire FA_cout_3163;
  wire FA_cout_3164;
  wire FA_cout_3165;
  wire FA_cout_3166;
  wire FA_cout_3167;
  wire FA_cout_3168;
  wire FA_cout_3169;
  wire FA_cout_3170;
  wire FA_cout_3171;
  wire FA_cout_3172;
  wire FA_cout_3173;
  wire FA_cout_3174;
  wire FA_cout_3175;
  wire FA_cout_3176;
  wire FA_cout_3177;
  wire FA_cout_3178;
  wire FA_cout_3179;
  wire FA_cout_3180;
  wire FA_cout_3181;
  wire FA_cout_3182;
  wire FA_cout_3183;
  wire FA_cout_3184;
  wire FA_cout_3185;
  wire FA_cout_3186;
  wire FA_cout_3187;
  wire FA_cout_3188;
  wire FA_cout_3189;
  wire FA_cout_3190;
  wire FA_cout_3191;
  wire FA_cout_3192;
  wire FA_cout_3193;
  wire FA_cout_3194;
  wire FA_cout_3195;
  wire FA_cout_3196;
  wire FA_cout_3197;
  wire FA_cout_3198;
  wire FA_cout_3199;
  wire FA_cout_3200;
  wire FA_cout_3201;
  wire FA_cout_3202;
  wire FA_cout_3203;
  wire FA_cout_3204;
  wire FA_cout_3205;
  wire FA_cout_3206;
  wire FA_cout_3207;
  wire FA_cout_3208;
  wire FA_cout_3209;
  wire FA_cout_3210;
  wire FA_cout_3211;
  wire FA_cout_3212;
  wire FA_cout_3213;
  wire FA_cout_3214;
  wire FA_cout_3215;
  wire FA_cout_3216;
  wire FA_cout_3217;
  wire FA_cout_3218;
  wire FA_cout_3219;
  wire FA_cout_3220;
  wire FA_cout_3221;
  wire FA_cout_3222;
  wire FA_cout_3223;
  wire FA_cout_3224;
  wire FA_cout_3225;
  wire FA_cout_3226;
  wire FA_cout_3227;
  wire FA_cout_3228;
  wire FA_cout_3229;
  wire FA_cout_3230;
  wire FA_cout_3231;
  wire FA_cout_3232;
  wire FA_cout_3233;
  wire FA_cout_3234;
  wire FA_cout_3235;
  wire FA_cout_3236;
  wire FA_cout_3237;
  wire FA_cout_3238;
  wire FA_cout_3239;
  wire FA_cout_3240;
  wire FA_cout_3241;
  wire FA_cout_3242;
  wire FA_cout_3243;
  wire FA_cout_3244;
  wire FA_cout_3245;
  wire FA_cout_3246;
  wire FA_cout_3247;
  wire FA_cout_3248;
  wire FA_cout_3249;
  wire FA_cout_3250;
  wire FA_cout_3251;
  wire FA_cout_3252;
  wire FA_cout_3253;
  wire FA_cout_3254;
  wire FA_cout_3255;
  wire FA_cout_3256;
  wire FA_cout_3257;
  wire FA_cout_3258;
  wire FA_cout_3259;
  wire FA_cout_3260;
  wire FA_cout_3261;
  wire FA_cout_3262;
  wire FA_cout_3263;
  wire FA_cout_3264;
  wire FA_cout_3265;
  wire FA_cout_3266;
  wire FA_cout_3267;
  wire FA_cout_3268;
  wire FA_cout_3269;
  wire FA_cout_3270;
  wire FA_cout_3271;
  wire FA_cout_3272;
  wire FA_cout_3273;
  wire FA_cout_3274;
  wire FA_cout_3275;
  wire FA_cout_3276;
  wire FA_cout_3277;
  wire FA_cout_3278;
  wire FA_cout_3279;
  wire FA_cout_3280;
  wire FA_cout_3281;
  wire FA_cout_3282;
  wire FA_cout_3283;
  wire FA_cout_3284;
  wire FA_cout_3285;
  wire FA_cout_3286;
  wire FA_cout_3287;
  wire FA_cout_3288;
  wire FA_cout_3289;
  wire FA_cout_3290;
  wire FA_cout_3291;
  wire FA_cout_3292;
  wire FA_cout_3293;
  wire FA_cout_3294;
  wire FA_cout_3295;
  wire FA_cout_3296;
  wire FA_cout_3297;
  wire FA_cout_3298;
  wire FA_cout_3299;
  wire FA_cout_3300;
  wire FA_cout_3301;
  wire FA_cout_3302;
  wire FA_cout_3303;
  wire FA_cout_3304;
  wire FA_cout_3305;
  wire FA_cout_3306;
  wire FA_cout_3307;
  wire FA_cout_3308;
  wire FA_cout_3309;
  wire FA_cout_3310;
  wire FA_cout_3311;
  wire FA_cout_3312;
  wire FA_cout_3313;
  wire FA_cout_3314;
  wire FA_cout_3315;
  wire FA_cout_3316;
  wire FA_cout_3317;
  wire FA_cout_3318;
  wire FA_cout_3319;
  wire FA_cout_3320;
  wire FA_cout_3321;
  wire FA_cout_3322;
  wire FA_cout_3323;
  wire FA_cout_3324;
  wire FA_cout_3325;
  wire FA_cout_3326;
  wire FA_cout_3327;
  wire FA_cout_3328;
  wire FA_cout_3329;
  wire FA_cout_3330;
  wire FA_cout_3331;
  wire FA_cout_3332;
  wire FA_cout_3333;
  wire FA_cout_3334;
  wire FA_cout_3335;
  wire FA_cout_3336;
  wire FA_cout_3337;
  wire FA_cout_3338;
  wire FA_cout_3339;
  wire FA_cout_3340;
  wire FA_cout_3341;
  wire FA_cout_3342;
  wire FA_cout_3343;
  wire FA_cout_3344;
  wire FA_cout_3345;
  wire FA_cout_3346;
  wire FA_cout_3347;
  wire FA_cout_3348;
  wire FA_cout_3349;
  wire FA_cout_3350;
  wire FA_cout_3351;
  wire FA_cout_3352;
  wire FA_cout_3353;
  wire FA_cout_3354;
  wire FA_cout_3355;
  wire FA_cout_3356;
  wire FA_cout_3357;
  wire FA_cout_3358;
  wire FA_cout_3359;
  wire FA_cout_3360;
  wire FA_cout_3361;
  wire FA_cout_3362;
  wire FA_cout_3363;
  wire FA_cout_3364;
  wire FA_cout_3365;
  wire FA_cout_3366;
  wire FA_cout_3367;
  wire FA_cout_3368;
  wire FA_cout_3369;
  wire FA_cout_3370;
  wire FA_cout_3371;
  wire FA_cout_3372;
  wire FA_cout_3373;
  wire FA_cout_3374;
  wire FA_cout_3375;
  wire FA_cout_3376;
  wire FA_cout_3377;
  wire FA_cout_3378;
  wire FA_cout_3379;
  wire FA_cout_3380;
  wire FA_cout_3381;
  wire FA_cout_3382;
  wire FA_cout_3383;
  wire FA_cout_3384;
  wire FA_cout_3385;
  wire FA_cout_3386;
  wire FA_cout_3387;
  wire FA_cout_3388;
  wire FA_cout_3389;
  wire FA_cout_3390;
  wire FA_cout_3391;
  wire FA_cout_3392;
  wire FA_cout_3393;
  wire FA_cout_3394;
  wire FA_cout_3395;
  wire FA_cout_3396;
  wire FA_cout_3397;
  wire FA_cout_3398;
  wire FA_cout_3399;
  wire FA_cout_3400;
  wire FA_cout_3401;
  wire FA_cout_3402;
  wire FA_cout_3403;
  wire FA_cout_3404;
  wire FA_cout_3405;
  wire FA_cout_3406;
  wire FA_cout_3407;
  wire FA_cout_3408;
  wire FA_cout_3409;
  wire FA_cout_3410;
  wire FA_cout_3411;
  wire FA_cout_3412;
  wire FA_cout_3413;
  wire FA_cout_3414;
  wire FA_cout_3415;
  wire FA_cout_3416;
  wire FA_cout_3417;
  wire FA_cout_3418;
  wire FA_cout_3419;
  wire FA_cout_3420;
  wire FA_cout_3421;
  wire FA_cout_3422;
  wire FA_cout_3423;
  wire FA_cout_3424;
  wire FA_cout_3425;
  wire FA_cout_3426;
  wire FA_cout_3427;
  wire FA_cout_3428;
  wire FA_cout_3429;
  wire FA_cout_3430;
  wire FA_cout_3431;
  wire FA_cout_3432;
  wire FA_cout_3433;
  wire FA_cout_3434;
  wire FA_cout_3435;
  wire FA_cout_3436;
  wire FA_cout_3437;
  wire FA_cout_3438;
  wire FA_cout_3439;
  wire FA_cout_3440;
  wire FA_cout_3441;
  wire FA_cout_3442;
  wire FA_cout_3443;
  wire FA_cout_3444;
  wire FA_cout_3445;
  wire FA_cout_3446;
  wire FA_cout_3447;
  wire FA_cout_3448;
  wire FA_cout_3449;
  wire FA_cout_3450;
  wire FA_cout_3451;
  wire FA_cout_3452;
  wire FA_cout_3453;
  wire FA_cout_3454;
  wire FA_cout_3455;
  wire FA_cout_3456;
  wire FA_cout_3457;
  wire FA_cout_3458;
  wire FA_cout_3459;
  wire FA_cout_3460;
  wire FA_cout_3461;
  wire FA_cout_3462;
  wire FA_cout_3463;
  wire FA_cout_3464;
  wire FA_cout_3465;
  wire FA_cout_3466;
  wire FA_cout_3467;
  wire FA_cout_3468;
  wire FA_cout_3469;
  wire FA_cout_3470;
  wire FA_cout_3471;
  wire FA_cout_3472;
  wire FA_cout_3473;
  wire FA_cout_3474;
  wire FA_cout_3475;
  wire FA_cout_3476;
  wire FA_cout_3477;
  wire FA_cout_3478;
  wire FA_cout_3479;
  wire FA_cout_3480;
  wire FA_cout_3481;
  wire FA_cout_3482;
  wire FA_cout_3483;
  wire FA_cout_3484;
  wire FA_cout_3485;
  wire FA_cout_3486;
  wire FA_cout_3487;
  wire FA_cout_3488;
  wire FA_cout_3489;
  wire FA_cout_3490;
  wire FA_cout_3491;
  wire FA_cout_3492;
  wire FA_cout_3493;
  wire FA_cout_3494;
  wire FA_cout_3495;
  wire FA_cout_3496;
  wire FA_cout_3497;
  wire FA_cout_3498;
  wire FA_cout_3499;
  wire FA_cout_3500;
  wire FA_cout_3501;
  wire FA_cout_3502;
  wire FA_cout_3503;
  wire FA_cout_3504;
  wire FA_cout_3505;
  wire FA_cout_3506;
  wire FA_cout_3507;
  wire FA_cout_3508;
  wire FA_cout_3509;
  wire FA_cout_3510;
  wire FA_cout_3511;
  wire FA_cout_3512;
  wire FA_cout_3513;
  wire FA_cout_3514;
  wire FA_cout_3515;
  wire FA_cout_3516;
  wire FA_cout_3517;
  wire FA_cout_3518;
  wire FA_cout_3519;
  wire FA_cout_3520;
  wire FA_cout_3521;
  wire FA_cout_3522;
  wire FA_cout_3523;
  wire FA_cout_3524;
  wire FA_cout_3525;
  wire FA_cout_3526;
  wire FA_cout_3527;
  wire FA_cout_3528;
  wire FA_cout_3529;
  wire FA_cout_3530;
  wire FA_cout_3531;
  wire FA_cout_3532;
  wire FA_cout_3533;
  wire FA_cout_3534;
  wire FA_cout_3535;
  wire FA_cout_3536;
  wire FA_cout_3537;
  wire FA_cout_3538;
  wire FA_cout_3539;
  wire FA_cout_3540;
  wire FA_cout_3541;
  wire FA_cout_3542;
  wire FA_cout_3543;
  wire FA_cout_3544;
  wire FA_cout_3545;
  wire FA_cout_3546;
  wire FA_cout_3547;
  wire FA_cout_3548;
  wire FA_cout_3549;
  wire FA_cout_3550;
  wire FA_cout_3551;
  wire FA_cout_3552;
  wire FA_cout_3553;
  wire FA_cout_3554;
  wire FA_cout_3555;
  wire FA_cout_3556;
  wire FA_cout_3557;
  wire FA_cout_3558;
  wire FA_cout_3559;
  wire FA_cout_3560;
  wire FA_cout_3561;
  wire FA_cout_3562;
  wire FA_cout_3563;
  wire FA_cout_3564;
  wire FA_cout_3565;
  wire FA_cout_3566;
  wire FA_cout_3567;
  wire FA_cout_3568;
  wire FA_cout_3569;
  wire FA_cout_3570;
  wire FA_cout_3571;
  wire FA_cout_3572;
  wire FA_cout_3573;
  wire FA_cout_3574;
  wire FA_cout_3575;
  wire FA_cout_3576;
  wire FA_cout_3577;
  wire FA_cout_3578;
  wire FA_cout_3579;
  wire FA_cout_3580;
  wire FA_cout_3581;
  wire FA_cout_3582;
  wire FA_cout_3583;
  wire FA_cout_3584;
  wire FA_cout_3585;
  wire FA_cout_3586;
  wire FA_cout_3587;
  wire FA_cout_3588;
  wire FA_cout_3589;
  wire FA_cout_3590;
  wire FA_cout_3591;
  wire FA_cout_3592;
  wire FA_cout_3593;
  wire FA_cout_3594;
  wire FA_cout_3595;
  wire FA_cout_3596;
  wire FA_cout_3597;
  wire FA_cout_3598;
  wire FA_cout_3599;
  wire FA_cout_3600;
  wire FA_cout_3601;
  wire FA_cout_3602;
  wire FA_cout_3603;
  wire FA_cout_3604;
  wire FA_cout_3605;
  wire FA_cout_3606;
  wire FA_cout_3607;
  wire FA_cout_3608;
  wire FA_cout_3609;
  wire FA_cout_3610;
  wire FA_cout_3611;
  wire FA_cout_3612;
  wire FA_cout_3613;
  wire FA_cout_3614;
  wire FA_cout_3615;
  wire FA_cout_3616;
  wire FA_cout_3617;
  wire FA_cout_3618;
  wire FA_cout_3619;
  wire FA_cout_3620;
  wire FA_cout_3621;
  wire FA_cout_3622;
  wire FA_cout_3623;
  wire FA_cout_3624;
  wire FA_cout_3625;
  wire FA_cout_3626;
  wire FA_cout_3627;
  wire FA_cout_3628;
  wire FA_cout_3629;
  wire FA_cout_3630;
  wire FA_cout_3631;
  wire FA_cout_3632;
  wire FA_cout_3633;
  wire FA_cout_3634;
  wire FA_cout_3635;
  wire FA_cout_3636;
  wire FA_cout_3637;
  wire FA_cout_3638;
  wire FA_cout_3639;
  wire FA_cout_3640;
  wire FA_cout_3641;
  wire FA_cout_3642;
  wire FA_cout_3643;
  wire FA_cout_3644;
  wire FA_cout_3645;
  wire FA_cout_3646;
  wire FA_cout_3647;
  wire FA_cout_3648;
  wire FA_cout_3649;
  wire FA_cout_3650;
  wire FA_cout_3651;
  wire FA_cout_3652;
  wire FA_cout_3653;
  wire FA_cout_3654;
  wire FA_cout_3655;
  wire FA_cout_3656;
  wire FA_cout_3657;
  wire FA_cout_3658;
  wire FA_cout_3659;
  wire FA_cout_3660;
  wire FA_cout_3661;
  wire FA_cout_3662;
  wire FA_cout_3663;
  wire FA_cout_3664;
  wire FA_cout_3665;
  wire FA_cout_3666;
  wire FA_cout_3667;
  wire FA_cout_3668;
  wire FA_cout_3669;
  wire FA_cout_3670;
  wire FA_cout_3671;
  wire FA_cout_3672;
  wire FA_cout_3673;
  wire FA_cout_3674;
  wire FA_cout_3675;
  wire FA_cout_3676;
  wire FA_cout_3677;
  wire FA_cout_3678;
  wire FA_cout_3679;
  wire FA_cout_3680;
  wire FA_cout_3681;
  wire FA_cout_3682;
  wire FA_cout_3683;
  wire FA_cout_3684;
  wire FA_cout_3685;
  wire FA_cout_3686;
  wire FA_cout_3687;
  wire FA_cout_3688;
  wire FA_cout_3689;
  wire FA_cout_3690;
  wire FA_cout_3691;
  wire FA_cout_3692;
  wire FA_cout_3693;
  wire FA_cout_3694;
  wire FA_cout_3695;
  wire FA_cout_3696;
  wire FA_cout_3697;
  wire FA_cout_3698;
  wire FA_cout_3699;
  wire FA_cout_3700;
  wire FA_cout_3701;
  wire FA_cout_3702;
  wire FA_cout_3703;
  wire FA_cout_3704;
  wire FA_cout_3705;
  wire FA_cout_3706;
  wire FA_cout_3707;
  wire FA_cout_3708;
  wire FA_cout_3709;
  wire FA_cout_3710;
  wire FA_cout_3711;
  wire FA_cout_3712;
  wire FA_cout_3713;
  wire FA_cout_3714;
  wire FA_cout_3715;
  wire FA_cout_3716;
  wire FA_cout_3717;
  wire FA_cout_3718;
  wire FA_cout_3719;
  wire FA_cout_3720;
  wire FA_cout_3721;
  wire FA_cout_3722;
  wire FA_cout_3723;
  wire FA_cout_3724;
  wire FA_cout_3725;
  wire FA_cout_3726;
  wire FA_cout_3727;
  wire FA_cout_3728;
  wire FA_cout_3729;
  wire FA_cout_3730;
  wire FA_cout_3731;
  wire FA_cout_3732;
  wire FA_cout_3733;
  wire FA_cout_3734;
  wire FA_cout_3735;
  wire FA_cout_3736;
  wire FA_cout_3737;
  wire FA_cout_3738;
  wire FA_cout_3739;
  wire FA_cout_3740;
  wire FA_cout_3741;
  wire FA_cout_3742;
  wire FA_cout_3743;
  wire FA_cout_3744;
  wire FA_cout_3745;
  wire FA_cout_3746;
  wire FA_cout_3747;
  wire FA_cout_3748;
  wire FA_cout_3749;
  wire FA_cout_3750;
  wire FA_cout_3751;
  wire FA_cout_3752;
  wire FA_cout_3753;
  wire FA_cout_3754;
  wire FA_cout_3755;
  wire FA_cout_3756;
  wire FA_cout_3757;
  wire FA_cout_3758;
  wire FA_cout_3759;
  wire FA_cout_3760;
  wire FA_cout_3761;
  wire FA_cout_3762;
  wire FA_cout_3763;
  wire FA_cout_3764;
  wire FA_cout_3765;
  wire FA_cout_3766;
  wire FA_cout_3767;
  wire FA_cout_3768;
  wire FA_cout_3769;
  wire FA_cout_3770;
  wire FA_cout_3771;
  wire FA_cout_3772;
  wire FA_cout_3773;
  wire FA_cout_3774;
  wire FA_cout_3775;
  wire FA_cout_3776;
  wire FA_cout_3777;
  wire FA_cout_3778;
  wire FA_cout_3779;
  wire FA_cout_3780;
  wire FA_cout_3781;
  wire FA_cout_3782;
  wire FA_cout_3783;
  wire FA_cout_3784;
  wire FA_cout_3785;
  wire FA_cout_3786;
  wire FA_cout_3787;
  wire FA_cout_3788;
  wire FA_cout_3789;
  wire FA_cout_3790;
  wire FA_cout_3791;
  wire FA_cout_3792;
  wire FA_cout_3793;
  wire FA_cout_3794;
  wire FA_cout_3795;
  wire FA_cout_3796;
  wire FA_cout_3797;
  wire FA_cout_3798;
  wire FA_cout_3799;
  wire FA_cout_3800;
  wire FA_cout_3801;
  wire FA_cout_3802;
  wire FA_cout_3803;
  wire FA_cout_3804;
  wire FA_cout_3805;
  wire FA_cout_3806;
  wire FA_cout_3807;
  wire FA_cout_3808;
  wire FA_cout_3809;
  wire FA_cout_3810;
  wire FA_cout_3811;
  wire FA_cout_3812;
  wire FA_cout_3813;
  wire FA_cout_3814;
  wire FA_cout_3815;
  wire FA_cout_3816;
  wire FA_cout_3817;
  wire FA_cout_3818;
  wire FA_cout_3819;
  wire FA_cout_3820;
  wire FA_cout_3821;
  wire FA_cout_3822;
  wire FA_cout_3823;
  wire FA_cout_3824;
  wire FA_cout_3825;
  wire FA_cout_3826;
  wire FA_cout_3827;
  wire FA_cout_3828;
  wire FA_cout_3829;
  wire FA_cout_3830;
  wire FA_cout_3831;
  wire FA_cout_3832;
  wire FA_cout_3833;
  wire FA_cout_3834;
  wire FA_cout_3835;
  wire FA_cout_3836;
  wire FA_cout_3837;
  wire FA_cout_3838;
  wire FA_cout_3839;
  wire FA_cout_3840;
  wire FA_cout_3841;
  wire FA_cout_3842;
  wire FA_cout_3843;
  wire HA_out_0;
  wire HA_out_1;
  wire HA_out_2;
  wire HA_out_3;
  wire HA_out_4;
  wire HA_out_5;
  wire HA_out_6;
  wire HA_out_7;
  wire HA_out_8;
  wire HA_out_9;
  wire HA_out_10;
  wire HA_out_11;
  wire HA_out_12;
  wire HA_out_13;
  wire HA_out_14;
  wire HA_out_15;
  wire HA_out_16;
  wire HA_out_17;
  wire HA_out_18;
  wire HA_out_19;
  wire HA_out_20;
  wire HA_out_21;
  wire HA_out_22;
  wire HA_out_23;
  wire HA_out_24;
  wire HA_out_25;
  wire HA_out_26;
  wire HA_out_27;
  wire HA_out_28;
  wire HA_out_29;
  wire HA_out_30;
  wire HA_out_31;
  wire HA_out_32;
  wire HA_out_33;
  wire HA_out_34;
  wire HA_out_35;
  wire HA_out_36;
  wire HA_out_37;
  wire HA_out_38;
  wire HA_out_39;
  wire HA_out_40;
  wire HA_out_41;
  wire HA_out_42;
  wire HA_out_43;
  wire HA_out_44;
  wire HA_out_45;
  wire HA_out_46;
  wire HA_out_47;
  wire HA_out_48;
  wire HA_out_49;
  wire HA_out_50;
  wire HA_out_51;
  wire HA_out_52;
  wire HA_out_53;
  wire HA_out_54;
  wire HA_out_55;
  wire HA_out_56;
  wire HA_out_57;
  wire HA_out_58;
  wire HA_out_59;
  wire HA_out_60;
  wire HA_out_61;
  wire HA_out_62;
  wire HA_out_63;
  wire HA_out_64;
  wire HA_out_65;
  wire HA_out_66;
  wire HA_out_67;
  wire HA_out_68;
  wire HA_out_69;
  wire HA_out_70;
  wire HA_out_71;
  wire HA_out_72;
  wire HA_out_73;
  wire HA_out_74;
  wire HA_out_75;
  wire HA_out_76;
  wire HA_out_77;
  wire HA_out_78;
  wire HA_out_79;
  wire HA_out_80;
  wire HA_out_81;
  wire HA_out_82;
  wire HA_out_83;
  wire HA_out_84;
  wire HA_out_85;
  wire HA_out_86;
  wire HA_out_87;
  wire HA_out_88;
  wire HA_out_89;
  wire HA_out_90;
  wire HA_out_91;
  wire HA_out_92;
  wire HA_out_93;
  wire HA_out_94;
  wire HA_out_95;
  wire HA_out_96;
  wire HA_out_97;
  wire HA_out_98;
  wire HA_out_99;
  wire HA_out_100;
  wire HA_out_101;
  wire HA_out_102;
  wire HA_out_103;
  wire HA_out_104;
  wire HA_out_105;
  wire HA_out_106;
  wire HA_out_107;
  wire HA_out_108;
  wire HA_out_109;
  wire HA_out_110;
  wire HA_out_111;
  wire HA_out_112;
  wire HA_out_113;
  wire HA_out_114;
  wire HA_out_115;
  wire HA_out_116;
  wire HA_out_117;
  wire HA_out_118;
  wire HA_out_119;
  wire HA_out_120;
  wire HA_out_121;
  wire HA_out_122;
  wire HA_out_123;
  wire HA_out_124;
  wire HA_out_125;
  wire HA_out_126;
  wire HA_out_127;
  wire HA_out_128;
  wire HA_out_129;
  wire HA_out_130;
  wire HA_out_131;
  wire HA_out_132;
  wire HA_out_133;
  wire HA_out_134;
  wire HA_out_135;
  wire HA_out_136;
  wire HA_out_137;
  wire HA_out_138;
  wire HA_out_139;
  wire HA_out_140;
  wire HA_out_141;
  wire HA_out_142;
  wire HA_out_143;
  wire HA_out_144;
  wire HA_out_145;
  wire HA_out_146;
  wire HA_out_147;
  wire HA_out_148;
  wire HA_out_149;
  wire HA_out_150;
  wire HA_out_151;
  wire HA_out_152;
  wire HA_out_153;
  wire HA_out_154;
  wire HA_out_155;
  wire HA_out_156;
  wire HA_out_157;
  wire HA_out_158;
  wire HA_out_159;
  wire HA_out_160;
  wire HA_out_161;
  wire HA_out_162;
  wire HA_out_163;
  wire HA_out_164;
  wire HA_out_165;
  wire HA_out_166;
  wire HA_out_167;
  wire HA_out_168;
  wire HA_out_169;
  wire HA_out_170;
  wire HA_out_171;
  wire HA_out_172;
  wire HA_out_173;
  wire HA_out_174;
  wire HA_out_175;
  wire HA_out_176;
  wire HA_out_177;
  wire HA_out_178;
  wire HA_out_179;
  wire HA_out_180;
  wire HA_out_181;
  wire HA_out_182;
  wire HA_out_183;
  wire HA_out_184;
  wire HA_out_185;
  wire HA_out_186;
  wire HA_out_187;
  wire HA_out_188;
  wire HA_out_189;
  wire HA_out_190;
  wire HA_out_191;
  wire HA_out_192;
  wire HA_out_193;
  wire HA_out_194;
  wire HA_out_195;
  wire HA_out_196;
  wire HA_out_197;
  wire HA_out_198;
  wire HA_out_199;
  wire HA_out_200;
  wire HA_out_201;
  wire HA_out_202;
  wire HA_out_203;
  wire HA_out_204;
  wire HA_out_205;
  wire HA_out_206;
  wire HA_out_207;
  wire HA_out_208;
  wire HA_out_209;
  wire HA_out_210;
  wire HA_out_211;
  wire HA_out_212;
  wire HA_out_213;
  wire HA_out_214;
  wire HA_out_215;
  wire HA_out_216;
  wire HA_out_217;
  wire HA_out_218;
  wire HA_out_219;
  wire HA_out_220;
  wire HA_out_221;
  wire HA_out_222;
  wire HA_out_223;
  wire HA_out_224;
  wire HA_out_225;
  wire HA_out_226;
  wire HA_out_227;
  wire HA_out_228;
  wire HA_out_229;
  wire HA_out_230;
  wire HA_out_231;
  wire HA_out_232;
  wire HA_out_233;
  wire HA_out_234;
  wire HA_out_235;
  wire HA_out_236;
  wire HA_out_237;
  wire HA_out_238;
  wire HA_out_239;
  wire HA_out_240;
  wire HA_out_241;
  wire HA_out_242;
  wire HA_out_243;
  wire HA_out_244;
  wire HA_out_245;
  wire HA_out_246;
  wire HA_out_247;
  wire HA_out_248;
  wire HA_out_249;
  wire HA_out_250;
  wire HA_out_251;
  wire HA_out_252;
  wire HA_out_253;
  wire HA_out_254;
  wire HA_out_255;
  wire HA_out_256;
  wire HA_out_257;
  wire HA_out_258;
  wire HA_out_259;
  wire HA_out_260;
  wire HA_out_261;
  wire HA_out_262;
  wire HA_out_263;
  wire HA_out_264;
  wire HA_out_265;
  wire HA_out_266;
  wire HA_out_267;
  wire HA_out_268;
  wire HA_out_269;
  wire HA_out_270;
  wire HA_out_271;
  wire HA_out_272;
  wire HA_out_273;
  wire HA_out_274;
  wire HA_out_275;
  wire HA_out_276;
  wire HA_out_277;
  wire HA_out_278;
  wire HA_out_279;
  wire HA_out_280;
  wire HA_out_281;
  wire HA_out_282;
  wire HA_out_283;
  wire HA_out_284;
  wire HA_out_285;
  wire HA_out_286;
  wire HA_out_287;
  wire HA_out_288;
  wire HA_out_289;
  wire HA_out_290;
  wire HA_out_291;
  wire HA_out_292;
  wire HA_out_293;
  wire HA_out_294;
  wire HA_out_295;
  wire HA_out_296;
  wire HA_out_297;
  wire HA_out_298;
  wire HA_out_299;
  wire HA_out_300;
  wire HA_out_301;
  wire HA_out_302;
  wire HA_out_303;
  wire HA_out_304;
  wire HA_out_305;
  wire HA_out_306;
  wire HA_out_307;
  wire HA_out_308;
  wire HA_out_309;
  wire HA_out_310;
  wire HA_out_311;
  wire HA_out_312;
  wire HA_out_313;
  wire HA_out_314;
  wire HA_out_315;
  wire HA_out_316;
  wire HA_out_317;
  wire HA_out_318;
  wire HA_out_319;
  wire HA_out_320;
  wire HA_out_321;
  wire HA_out_322;
  wire HA_out_323;
  wire HA_out_324;
  wire HA_out_325;
  wire HA_out_326;
  wire HA_out_327;
  wire HA_out_328;
  wire HA_out_329;
  wire HA_out_330;
  wire HA_out_331;
  wire HA_out_332;
  wire HA_out_333;
  wire HA_out_334;
  wire HA_out_335;
  wire HA_out_336;
  wire HA_out_337;
  wire HA_out_338;
  wire HA_out_339;
  wire HA_out_340;
  wire HA_out_341;
  wire HA_out_342;
  wire HA_out_343;
  wire HA_out_344;
  wire HA_out_345;
  wire HA_out_346;
  wire HA_out_347;
  wire HA_out_348;
  wire HA_out_349;
  wire HA_out_350;
  wire HA_out_351;
  wire HA_out_352;
  wire HA_out_353;
  wire HA_out_354;
  wire HA_out_355;
  wire HA_out_356;
  wire HA_out_357;
  wire HA_out_358;
  wire HA_out_359;
  wire HA_out_360;
  wire HA_out_361;
  wire HA_out_362;
  wire HA_out_363;
  wire HA_out_364;
  wire HA_out_365;
  wire HA_out_366;
  wire HA_out_367;
  wire HA_out_368;
  wire HA_out_369;
  wire HA_out_370;
  wire HA_out_371;
  wire HA_out_372;
  wire HA_out_373;
  wire HA_out_374;
  wire HA_out_375;
  wire HA_out_376;
  wire HA_out_377;
  wire HA_out_378;
  wire HA_out_379;
  wire HA_out_380;
  wire HA_out_381;
  wire HA_out_382;
  wire HA_out_383;
  wire HA_out_384;
  wire HA_out_385;
  wire HA_out_386;
  wire HA_out_387;
  wire HA_out_388;
  wire HA_out_389;
  wire HA_out_390;
  wire HA_out_391;
  wire HA_out_392;
  wire HA_out_393;
  wire HA_out_394;
  wire HA_out_395;
  wire HA_out_396;
  wire HA_out_397;
  wire HA_out_398;
  wire HA_out_399;
  wire HA_out_400;
  wire HA_out_401;
  wire HA_out_402;
  wire HA_out_403;
  wire HA_out_404;
  wire HA_out_405;
  wire HA_out_406;
  wire HA_out_407;
  wire HA_out_408;
  wire HA_out_409;
  wire HA_out_410;
  wire HA_out_411;
  wire HA_out_412;
  wire HA_out_413;
  wire HA_out_414;
  wire HA_out_415;
  wire HA_out_416;
  wire HA_out_417;
  wire HA_out_418;
  wire HA_out_419;
  wire HA_out_420;
  wire HA_out_421;
  wire HA_out_422;
  wire HA_out_423;
  wire HA_out_424;
  wire HA_out_425;
  wire HA_out_426;
  wire HA_out_427;
  wire HA_out_428;
  wire HA_out_429;
  wire HA_out_430;
  wire HA_out_431;
  wire HA_out_432;
  wire HA_out_433;
  wire HA_out_434;
  wire HA_out_435;
  wire HA_out_436;
  wire HA_out_437;
  wire HA_out_438;
  wire HA_out_439;
  wire HA_out_440;
  wire HA_out_441;
  wire HA_out_442;
  wire HA_out_443;
  wire HA_out_444;
  wire HA_out_445;
  wire HA_out_446;
  wire HA_out_447;
  wire HA_out_448;
  wire HA_out_449;
  wire HA_out_450;
  wire HA_out_451;
  wire HA_out_452;
  wire HA_out_453;
  wire HA_out_454;
  wire HA_out_455;
  wire HA_out_456;
  wire HA_out_457;
  wire HA_out_458;
  wire HA_out_459;
  wire HA_out_460;
  wire HA_out_461;
  wire HA_out_462;
  wire HA_out_463;
  wire HA_out_464;
  wire HA_out_465;
  wire HA_out_466;
  wire HA_out_467;
  wire HA_out_468;
  wire HA_out_469;
  wire HA_out_470;
  wire HA_out_471;
  wire HA_out_472;
  wire HA_out_473;
  wire HA_out_474;
  wire HA_out_475;
  wire HA_out_476;
  wire HA_out_477;
  wire HA_out_478;
  wire HA_out_479;
  wire HA_out_480;
  wire HA_out_481;
  wire HA_out_482;
  wire HA_out_483;
  wire HA_out_484;
  wire HA_out_485;
  wire HA_out_486;
  wire HA_out_487;
  wire HA_out_488;
  wire HA_out_489;
  wire HA_out_490;
  wire HA_out_491;
  wire HA_out_492;
  wire HA_out_493;
  wire HA_out_494;
  wire HA_out_495;
  wire HA_out_496;
  wire HA_out_497;
  wire HA_out_498;
  wire HA_out_499;
  wire HA_out_500;
  wire HA_out_501;
  wire HA_out_502;
  wire HA_out_503;
  wire HA_out_504;
  wire HA_out_505;
  wire HA_out_506;
  wire HA_out_507;
  wire HA_out_508;
  wire HA_out_509;
  wire HA_out_510;
  wire HA_out_511;
  wire HA_out_512;
  wire HA_out_513;
  wire HA_out_514;
  wire HA_out_515;
  wire HA_out_516;
  wire HA_out_517;
  wire HA_out_518;
  wire HA_out_519;
  wire HA_out_520;
  wire HA_out_521;
  wire HA_out_522;
  wire HA_out_523;
  wire HA_out_524;
  wire HA_out_525;
  wire HA_out_526;
  wire HA_out_527;
  wire HA_out_528;
  wire HA_out_529;
  wire HA_out_530;
  wire HA_out_531;
  wire HA_out_532;
  wire HA_out_533;
  wire HA_out_534;
  wire HA_out_535;
  wire HA_out_536;
  wire HA_out_537;
  wire HA_out_538;
  wire HA_out_539;
  wire HA_out_540;
  wire HA_out_541;
  wire HA_out_542;
  wire HA_out_543;
  wire HA_out_544;
  wire HA_out_545;
  wire HA_out_546;
  wire HA_out_547;
  wire HA_out_548;
  wire HA_out_549;
  wire HA_out_550;
  wire HA_out_551;
  wire HA_out_552;
  wire HA_out_553;
  wire HA_out_554;
  wire HA_out_555;
  wire HA_out_556;
  wire HA_out_557;
  wire HA_out_558;
  wire HA_out_559;
  wire HA_out_560;
  wire HA_cout_0;
  wire HA_cout_1;
  wire HA_cout_2;
  wire HA_cout_3;
  wire HA_cout_4;
  wire HA_cout_5;
  wire HA_cout_6;
  wire HA_cout_7;
  wire HA_cout_8;
  wire HA_cout_9;
  wire HA_cout_10;
  wire HA_cout_11;
  wire HA_cout_12;
  wire HA_cout_13;
  wire HA_cout_14;
  wire HA_cout_15;
  wire HA_cout_16;
  wire HA_cout_17;
  wire HA_cout_18;
  wire HA_cout_19;
  wire HA_cout_20;
  wire HA_cout_21;
  wire HA_cout_22;
  wire HA_cout_23;
  wire HA_cout_24;
  wire HA_cout_25;
  wire HA_cout_26;
  wire HA_cout_27;
  wire HA_cout_28;
  wire HA_cout_29;
  wire HA_cout_30;
  wire HA_cout_31;
  wire HA_cout_32;
  wire HA_cout_33;
  wire HA_cout_34;
  wire HA_cout_35;
  wire HA_cout_36;
  wire HA_cout_37;
  wire HA_cout_38;
  wire HA_cout_39;
  wire HA_cout_40;
  wire HA_cout_41;
  wire HA_cout_42;
  wire HA_cout_43;
  wire HA_cout_44;
  wire HA_cout_45;
  wire HA_cout_46;
  wire HA_cout_47;
  wire HA_cout_48;
  wire HA_cout_49;
  wire HA_cout_50;
  wire HA_cout_51;
  wire HA_cout_52;
  wire HA_cout_53;
  wire HA_cout_54;
  wire HA_cout_55;
  wire HA_cout_56;
  wire HA_cout_57;
  wire HA_cout_58;
  wire HA_cout_59;
  wire HA_cout_60;
  wire HA_cout_61;
  wire HA_cout_62;
  wire HA_cout_63;
  wire HA_cout_64;
  wire HA_cout_65;
  wire HA_cout_66;
  wire HA_cout_67;
  wire HA_cout_68;
  wire HA_cout_69;
  wire HA_cout_70;
  wire HA_cout_71;
  wire HA_cout_72;
  wire HA_cout_73;
  wire HA_cout_74;
  wire HA_cout_75;
  wire HA_cout_76;
  wire HA_cout_77;
  wire HA_cout_78;
  wire HA_cout_79;
  wire HA_cout_80;
  wire HA_cout_81;
  wire HA_cout_82;
  wire HA_cout_83;
  wire HA_cout_84;
  wire HA_cout_85;
  wire HA_cout_86;
  wire HA_cout_87;
  wire HA_cout_88;
  wire HA_cout_89;
  wire HA_cout_90;
  wire HA_cout_91;
  wire HA_cout_92;
  wire HA_cout_93;
  wire HA_cout_94;
  wire HA_cout_95;
  wire HA_cout_96;
  wire HA_cout_97;
  wire HA_cout_98;
  wire HA_cout_99;
  wire HA_cout_100;
  wire HA_cout_101;
  wire HA_cout_102;
  wire HA_cout_103;
  wire HA_cout_104;
  wire HA_cout_105;
  wire HA_cout_106;
  wire HA_cout_107;
  wire HA_cout_108;
  wire HA_cout_109;
  wire HA_cout_110;
  wire HA_cout_111;
  wire HA_cout_112;
  wire HA_cout_113;
  wire HA_cout_114;
  wire HA_cout_115;
  wire HA_cout_116;
  wire HA_cout_117;
  wire HA_cout_118;
  wire HA_cout_119;
  wire HA_cout_120;
  wire HA_cout_121;
  wire HA_cout_122;
  wire HA_cout_123;
  wire HA_cout_124;
  wire HA_cout_125;
  wire HA_cout_126;
  wire HA_cout_127;
  wire HA_cout_128;
  wire HA_cout_129;
  wire HA_cout_130;
  wire HA_cout_131;
  wire HA_cout_132;
  wire HA_cout_133;
  wire HA_cout_134;
  wire HA_cout_135;
  wire HA_cout_136;
  wire HA_cout_137;
  wire HA_cout_138;
  wire HA_cout_139;
  wire HA_cout_140;
  wire HA_cout_141;
  wire HA_cout_142;
  wire HA_cout_143;
  wire HA_cout_144;
  wire HA_cout_145;
  wire HA_cout_146;
  wire HA_cout_147;
  wire HA_cout_148;
  wire HA_cout_149;
  wire HA_cout_150;
  wire HA_cout_151;
  wire HA_cout_152;
  wire HA_cout_153;
  wire HA_cout_154;
  wire HA_cout_155;
  wire HA_cout_156;
  wire HA_cout_157;
  wire HA_cout_158;
  wire HA_cout_159;
  wire HA_cout_160;
  wire HA_cout_161;
  wire HA_cout_162;
  wire HA_cout_163;
  wire HA_cout_164;
  wire HA_cout_165;
  wire HA_cout_166;
  wire HA_cout_167;
  wire HA_cout_168;
  wire HA_cout_169;
  wire HA_cout_170;
  wire HA_cout_171;
  wire HA_cout_172;
  wire HA_cout_173;
  wire HA_cout_174;
  wire HA_cout_175;
  wire HA_cout_176;
  wire HA_cout_177;
  wire HA_cout_178;
  wire HA_cout_179;
  wire HA_cout_180;
  wire HA_cout_181;
  wire HA_cout_182;
  wire HA_cout_183;
  wire HA_cout_184;
  wire HA_cout_185;
  wire HA_cout_186;
  wire HA_cout_187;
  wire HA_cout_188;
  wire HA_cout_189;
  wire HA_cout_190;
  wire HA_cout_191;
  wire HA_cout_192;
  wire HA_cout_193;
  wire HA_cout_194;
  wire HA_cout_195;
  wire HA_cout_196;
  wire HA_cout_197;
  wire HA_cout_198;
  wire HA_cout_199;
  wire HA_cout_200;
  wire HA_cout_201;
  wire HA_cout_202;
  wire HA_cout_203;
  wire HA_cout_204;
  wire HA_cout_205;
  wire HA_cout_206;
  wire HA_cout_207;
  wire HA_cout_208;
  wire HA_cout_209;
  wire HA_cout_210;
  wire HA_cout_211;
  wire HA_cout_212;
  wire HA_cout_213;
  wire HA_cout_214;
  wire HA_cout_215;
  wire HA_cout_216;
  wire HA_cout_217;
  wire HA_cout_218;
  wire HA_cout_219;
  wire HA_cout_220;
  wire HA_cout_221;
  wire HA_cout_222;
  wire HA_cout_223;
  wire HA_cout_224;
  wire HA_cout_225;
  wire HA_cout_226;
  wire HA_cout_227;
  wire HA_cout_228;
  wire HA_cout_229;
  wire HA_cout_230;
  wire HA_cout_231;
  wire HA_cout_232;
  wire HA_cout_233;
  wire HA_cout_234;
  wire HA_cout_235;
  wire HA_cout_236;
  wire HA_cout_237;
  wire HA_cout_238;
  wire HA_cout_239;
  wire HA_cout_240;
  wire HA_cout_241;
  wire HA_cout_242;
  wire HA_cout_243;
  wire HA_cout_244;
  wire HA_cout_245;
  wire HA_cout_246;
  wire HA_cout_247;
  wire HA_cout_248;
  wire HA_cout_249;
  wire HA_cout_250;
  wire HA_cout_251;
  wire HA_cout_252;
  wire HA_cout_253;
  wire HA_cout_254;
  wire HA_cout_255;
  wire HA_cout_256;
  wire HA_cout_257;
  wire HA_cout_258;
  wire HA_cout_259;
  wire HA_cout_260;
  wire HA_cout_261;
  wire HA_cout_262;
  wire HA_cout_263;
  wire HA_cout_264;
  wire HA_cout_265;
  wire HA_cout_266;
  wire HA_cout_267;
  wire HA_cout_268;
  wire HA_cout_269;
  wire HA_cout_270;
  wire HA_cout_271;
  wire HA_cout_272;
  wire HA_cout_273;
  wire HA_cout_274;
  wire HA_cout_275;
  wire HA_cout_276;
  wire HA_cout_277;
  wire HA_cout_278;
  wire HA_cout_279;
  wire HA_cout_280;
  wire HA_cout_281;
  wire HA_cout_282;
  wire HA_cout_283;
  wire HA_cout_284;
  wire HA_cout_285;
  wire HA_cout_286;
  wire HA_cout_287;
  wire HA_cout_288;
  wire HA_cout_289;
  wire HA_cout_290;
  wire HA_cout_291;
  wire HA_cout_292;
  wire HA_cout_293;
  wire HA_cout_294;
  wire HA_cout_295;
  wire HA_cout_296;
  wire HA_cout_297;
  wire HA_cout_298;
  wire HA_cout_299;
  wire HA_cout_300;
  wire HA_cout_301;
  wire HA_cout_302;
  wire HA_cout_303;
  wire HA_cout_304;
  wire HA_cout_305;
  wire HA_cout_306;
  wire HA_cout_307;
  wire HA_cout_308;
  wire HA_cout_309;
  wire HA_cout_310;
  wire HA_cout_311;
  wire HA_cout_312;
  wire HA_cout_313;
  wire HA_cout_314;
  wire HA_cout_315;
  wire HA_cout_316;
  wire HA_cout_317;
  wire HA_cout_318;
  wire HA_cout_319;
  wire HA_cout_320;
  wire HA_cout_321;
  wire HA_cout_322;
  wire HA_cout_323;
  wire HA_cout_324;
  wire HA_cout_325;
  wire HA_cout_326;
  wire HA_cout_327;
  wire HA_cout_328;
  wire HA_cout_329;
  wire HA_cout_330;
  wire HA_cout_331;
  wire HA_cout_332;
  wire HA_cout_333;
  wire HA_cout_334;
  wire HA_cout_335;
  wire HA_cout_336;
  wire HA_cout_337;
  wire HA_cout_338;
  wire HA_cout_339;
  wire HA_cout_340;
  wire HA_cout_341;
  wire HA_cout_342;
  wire HA_cout_343;
  wire HA_cout_344;
  wire HA_cout_345;
  wire HA_cout_346;
  wire HA_cout_347;
  wire HA_cout_348;
  wire HA_cout_349;
  wire HA_cout_350;
  wire HA_cout_351;
  wire HA_cout_352;
  wire HA_cout_353;
  wire HA_cout_354;
  wire HA_cout_355;
  wire HA_cout_356;
  wire HA_cout_357;
  wire HA_cout_358;
  wire HA_cout_359;
  wire HA_cout_360;
  wire HA_cout_361;
  wire HA_cout_362;
  wire HA_cout_363;
  wire HA_cout_364;
  wire HA_cout_365;
  wire HA_cout_366;
  wire HA_cout_367;
  wire HA_cout_368;
  wire HA_cout_369;
  wire HA_cout_370;
  wire HA_cout_371;
  wire HA_cout_372;
  wire HA_cout_373;
  wire HA_cout_374;
  wire HA_cout_375;
  wire HA_cout_376;
  wire HA_cout_377;
  wire HA_cout_378;
  wire HA_cout_379;
  wire HA_cout_380;
  wire HA_cout_381;
  wire HA_cout_382;
  wire HA_cout_383;
  wire HA_cout_384;
  wire HA_cout_385;
  wire HA_cout_386;
  wire HA_cout_387;
  wire HA_cout_388;
  wire HA_cout_389;
  wire HA_cout_390;
  wire HA_cout_391;
  wire HA_cout_392;
  wire HA_cout_393;
  wire HA_cout_394;
  wire HA_cout_395;
  wire HA_cout_396;
  wire HA_cout_397;
  wire HA_cout_398;
  wire HA_cout_399;
  wire HA_cout_400;
  wire HA_cout_401;
  wire HA_cout_402;
  wire HA_cout_403;
  wire HA_cout_404;
  wire HA_cout_405;
  wire HA_cout_406;
  wire HA_cout_407;
  wire HA_cout_408;
  wire HA_cout_409;
  wire HA_cout_410;
  wire HA_cout_411;
  wire HA_cout_412;
  wire HA_cout_413;
  wire HA_cout_414;
  wire HA_cout_415;
  wire HA_cout_416;
  wire HA_cout_417;
  wire HA_cout_418;
  wire HA_cout_419;
  wire HA_cout_420;
  wire HA_cout_421;
  wire HA_cout_422;
  wire HA_cout_423;
  wire HA_cout_424;
  wire HA_cout_425;
  wire HA_cout_426;
  wire HA_cout_427;
  wire HA_cout_428;
  wire HA_cout_429;
  wire HA_cout_430;
  wire HA_cout_431;
  wire HA_cout_432;
  wire HA_cout_433;
  wire HA_cout_434;
  wire HA_cout_435;
  wire HA_cout_436;
  wire HA_cout_437;
  wire HA_cout_438;
  wire HA_cout_439;
  wire HA_cout_440;
  wire HA_cout_441;
  wire HA_cout_442;
  wire HA_cout_443;
  wire HA_cout_444;
  wire HA_cout_445;
  wire HA_cout_446;
  wire HA_cout_447;
  wire HA_cout_448;
  wire HA_cout_449;
  wire HA_cout_450;
  wire HA_cout_451;
  wire HA_cout_452;
  wire HA_cout_453;
  wire HA_cout_454;
  wire HA_cout_455;
  wire HA_cout_456;
  wire HA_cout_457;
  wire HA_cout_458;
  wire HA_cout_459;
  wire HA_cout_460;
  wire HA_cout_461;
  wire HA_cout_462;
  wire HA_cout_463;
  wire HA_cout_464;
  wire HA_cout_465;
  wire HA_cout_466;
  wire HA_cout_467;
  wire HA_cout_468;
  wire HA_cout_469;
  wire HA_cout_470;
  wire HA_cout_471;
  wire HA_cout_472;
  wire HA_cout_473;
  wire HA_cout_474;
  wire HA_cout_475;
  wire HA_cout_476;
  wire HA_cout_477;
  wire HA_cout_478;
  wire HA_cout_479;
  wire HA_cout_480;
  wire HA_cout_481;
  wire HA_cout_482;
  wire HA_cout_483;
  wire HA_cout_484;
  wire HA_cout_485;
  wire HA_cout_486;
  wire HA_cout_487;
  wire HA_cout_488;
  wire HA_cout_489;
  wire HA_cout_490;
  wire HA_cout_491;
  wire HA_cout_492;
  wire HA_cout_493;
  wire HA_cout_494;
  wire HA_cout_495;
  wire HA_cout_496;
  wire HA_cout_497;
  wire HA_cout_498;
  wire HA_cout_499;
  wire HA_cout_500;
  wire HA_cout_501;
  wire HA_cout_502;
  wire HA_cout_503;
  wire HA_cout_504;
  wire HA_cout_505;
  wire HA_cout_506;
  wire HA_cout_507;
  wire HA_cout_508;
  wire HA_cout_509;
  wire HA_cout_510;
  wire HA_cout_511;
  wire HA_cout_512;
  wire HA_cout_513;
  wire HA_cout_514;
  wire HA_cout_515;
  wire HA_cout_516;
  wire HA_cout_517;
  wire HA_cout_518;
  wire HA_cout_519;
  wire HA_cout_520;
  wire HA_cout_521;
  wire HA_cout_522;
  wire HA_cout_523;
  wire HA_cout_524;
  wire HA_cout_525;
  wire HA_cout_526;
  wire HA_cout_527;
  wire HA_cout_528;
  wire HA_cout_529;
  wire HA_cout_530;
  wire HA_cout_531;
  wire HA_cout_532;
  wire HA_cout_533;
  wire HA_cout_534;
  wire HA_cout_535;
  wire HA_cout_536;
  wire HA_cout_537;
  wire HA_cout_538;
  wire HA_cout_539;
  wire HA_cout_540;
  wire HA_cout_541;
  wire HA_cout_542;
  wire HA_cout_543;
  wire HA_cout_544;
  wire HA_cout_545;
  wire HA_cout_546;
  wire HA_cout_547;
  wire HA_cout_548;
  wire HA_cout_549;
  wire HA_cout_550;
  wire HA_cout_551;
  wire HA_cout_552;
  wire HA_cout_553;
  wire HA_cout_554;
  wire HA_cout_555;
  wire HA_cout_556;
  wire HA_cout_557;
  wire HA_cout_558;
  wire HA_cout_559;
  wire HA_cout_560;
  wire [64:0] inp_0;

  wire [64:0] inp_1;

  wire [64:0] inp_2;

  wire [64:0] inp_3;

  wire [64:0] inp_4;

  wire [64:0] inp_5;

  wire [64:0] inp_6;

  wire [64:0] inp_7;

  wire [64:0] inp_8;

  wire [64:0] inp_9;

  wire [64:0] inp_10;

  wire [64:0] inp_11;

  wire [64:0] inp_12;

  wire [64:0] inp_13;

  wire [64:0] inp_14;

  wire [64:0] inp_15;

  wire [64:0] inp_16;

  wire [64:0] inp_17;

  wire [64:0] inp_18;

  wire [64:0] inp_19;

  wire [64:0] inp_20;

  wire [64:0] inp_21;

  wire [64:0] inp_22;

  wire [64:0] inp_23;

  wire [64:0] inp_24;

  wire [64:0] inp_25;

  wire [64:0] inp_26;

  wire [64:0] inp_27;

  wire [64:0] inp_28;

  wire [64:0] inp_29;

  wire [64:0] inp_30;

  wire [64:0] inp_31;

  wire [64:0] inp_32;

  wire [64:0] inp_33;

  wire [64:0] inp_34;

  wire [64:0] inp_35;

  wire [64:0] inp_36;

  wire [64:0] inp_37;

  wire [64:0] inp_38;

  wire [64:0] inp_39;

  wire [64:0] inp_40;

  wire [64:0] inp_41;

  wire [64:0] inp_42;

  wire [64:0] inp_43;

  wire [64:0] inp_44;

  wire [64:0] inp_45;

  wire [64:0] inp_46;

  wire [64:0] inp_47;

  wire [64:0] inp_48;

  wire [64:0] inp_49;

  wire [64:0] inp_50;

  wire [64:0] inp_51;

  wire [64:0] inp_52;

  wire [64:0] inp_53;

  wire [64:0] inp_54;

  wire [64:0] inp_55;

  wire [64:0] inp_56;

  wire [64:0] inp_57;

  wire [64:0] inp_58;

  wire [64:0] inp_59;

  wire [64:0] inp_60;

  wire [64:0] inp_61;

  wire [64:0] inp_62;

  wire [64:0] inp_63;

  assign inp_0[51:0]=C[51:0] & {52{R[0]}};
  assign inp_0[52]=(C[52]|or1) && (R[0]);
  assign inp_0[63:53]=C[63:53] & {11{R[0]&and1}};
  assign inp_1[51:0]=C[51:0] & {52{R[1]}};
  assign inp_1[52]=(C[52]|or1) && (R[1]);
  assign inp_1[63:53]=C[63:53] & {11{R[1]&and1}};
  assign inp_2[51:0]=C[51:0] & {52{R[2]}};
  assign inp_2[52]=(C[52]|or1) && (R[2]);
  assign inp_2[63:53]=C[63:53] & {11{R[2]&and1}};
  assign inp_3[51:0]=C[51:0] & {52{R[3]}};
  assign inp_3[52]=(C[52]|or1) && (R[3]);
  assign inp_3[63:53]=C[63:53] & {11{R[3]&and1}};
  assign inp_4[51:0]=C[51:0] & {52{R[4]}};
  assign inp_4[52]=(C[52]|or1) && (R[4]);
  assign inp_4[63:53]=C[63:53] & {11{R[4]&and1}};
  assign inp_5[51:0]=C[51:0] & {52{R[5]}};
  assign inp_5[52]=(C[52]|or1) && (R[5]);
  assign inp_5[63:53]=C[63:53] & {11{R[5]&and1}};
  assign inp_6[51:0]=C[51:0] & {52{R[6]}};
  assign inp_6[52]=(C[52]|or1) && (R[6]);
  assign inp_6[63:53]=C[63:53] & {11{R[6]&and1}};
  assign inp_7[51:0]=C[51:0] & {52{R[7]}};
  assign inp_7[52]=(C[52]|or1) && (R[7]);
  assign inp_7[63:53]=C[63:53] & {11{R[7]&and1}};
  assign inp_8[51:0]=C[51:0] & {52{R[8]}};
  assign inp_8[52]=(C[52]|or1) && (R[8]);
  assign inp_8[63:53]=C[63:53] & {11{R[8]&and1}};
  assign inp_9[51:0]=C[51:0] & {52{R[9]}};
  assign inp_9[52]=(C[52]|or1) && (R[9]);
  assign inp_9[63:53]=C[63:53] & {11{R[9]&and1}};
  assign inp_10[51:0]=C[51:0] & {52{R[10]}};
  assign inp_10[52]=(C[52]|or1) && (R[10]);
  assign inp_10[63:53]=C[63:53] & {11{R[10]&and1}};
  assign inp_11[51:0]=C[51:0] & {52{R[11]}};
  assign inp_11[52]=(C[52]|or1) && (R[11]);
  assign inp_11[63:53]=C[63:53] & {11{R[11]&and1}};
  assign inp_12[51:0]=C[51:0] & {52{R[12]}};
  assign inp_12[52]=(C[52]|or1) && (R[12]);
  assign inp_12[63:53]=C[63:53] & {11{R[12]&and1}};
  assign inp_13[51:0]=C[51:0] & {52{R[13]}};
  assign inp_13[52]=(C[52]|or1) && (R[13]);
  assign inp_13[63:53]=C[63:53] & {11{R[13]&and1}};
  assign inp_14[51:0]=C[51:0] & {52{R[14]}};
  assign inp_14[52]=(C[52]|or1) && (R[14]);
  assign inp_14[63:53]=C[63:53] & {11{R[14]&and1}};
  assign inp_15[51:0]=C[51:0] & {52{R[15]}};
  assign inp_15[52]=(C[52]|or1) && (R[15]);
  assign inp_15[63:53]=C[63:53] & {11{R[15]&and1}};
  assign inp_16[51:0]=C[51:0] & {52{R[16]}};
  assign inp_16[52]=(C[52]|or1) && (R[16]);
  assign inp_16[63:53]=C[63:53] & {11{R[16]&and1}};
  assign inp_17[51:0]=C[51:0] & {52{R[17]}};
  assign inp_17[52]=(C[52]|or1) && (R[17]);
  assign inp_17[63:53]=C[63:53] & {11{R[17]&and1}};
  assign inp_18[51:0]=C[51:0] & {52{R[18]}};
  assign inp_18[52]=(C[52]|or1) && (R[18]);
  assign inp_18[63:53]=C[63:53] & {11{R[18]&and1}};
  assign inp_19[51:0]=C[51:0] & {52{R[19]}};
  assign inp_19[52]=(C[52]|or1) && (R[19]);
  assign inp_19[63:53]=C[63:53] & {11{R[19]&and1}};
  assign inp_20[51:0]=C[51:0] & {52{R[20]}};
  assign inp_20[52]=(C[52]|or1) && (R[20]);
  assign inp_20[63:53]=C[63:53] & {11{R[20]&and1}};
  assign inp_21[51:0]=C[51:0] & {52{R[21]}};
  assign inp_21[52]=(C[52]|or1) && (R[21]);
  assign inp_21[63:53]=C[63:53] & {11{R[21]&and1}};
  assign inp_22[51:0]=C[51:0] & {52{R[22]}};
  assign inp_22[52]=(C[52]|or1) && (R[22]);
  assign inp_22[63:53]=C[63:53] & {11{R[22]&and1}};
  assign inp_23[51:0]=C[51:0] & {52{R[23]}};
  assign inp_23[52]=(C[52]|or1) && (R[23]);
  assign inp_23[63:53]=C[63:53] & {11{R[23]&and1}};
  assign inp_24[51:0]=C[51:0] & {52{R[24]}};
  assign inp_24[52]=(C[52]|or1) && (R[24]);
  assign inp_24[63:53]=C[63:53] & {11{R[24]&and1}};
  assign inp_25[51:0]=C[51:0] & {52{R[25]}};
  assign inp_25[52]=(C[52]|or1) && (R[25]);
  assign inp_25[63:53]=C[63:53] & {11{R[25]&and1}};
  assign inp_26[51:0]=C[51:0] & {52{R[26]}};
  assign inp_26[52]=(C[52]|or1) && (R[26]);
  assign inp_26[63:53]=C[63:53] & {11{R[26]&and1}};
  assign inp_27[51:0]=C[51:0] & {52{R[27]}};
  assign inp_27[52]=(C[52]|or1) && (R[27]);
  assign inp_27[63:53]=C[63:53] & {11{R[27]&and1}};
  assign inp_28[51:0]=C[51:0] & {52{R[28]}};
  assign inp_28[52]=(C[52]|or1) && (R[28]);
  assign inp_28[63:53]=C[63:53] & {11{R[28]&and1}};
  assign inp_29[51:0]=C[51:0] & {52{R[29]}};
  assign inp_29[52]=(C[52]|or1) && (R[29]);
  assign inp_29[63:53]=C[63:53] & {11{R[29]&and1}};
  assign inp_30[51:0]=C[51:0] & {52{R[30]}};
  assign inp_30[52]=(C[52]|or1) && (R[30]);
  assign inp_30[63:53]=C[63:53] & {11{R[30]&and1}};
  assign inp_31[51:0]=C[51:0] & {52{R[31]}};
  assign inp_31[52]=(C[52]|or1) && (R[31]);
  assign inp_31[63:53]=C[63:53] & {11{R[31]&and1}};
  assign inp_32[51:0]=C[51:0] & {52{R[32]}};
  assign inp_32[52]=(C[52]|or1) && (R[32]);
  assign inp_32[63:53]=C[63:53] & {11{R[32]&and1}};
  assign inp_33[51:0]=C[51:0] & {52{R[33]}};
  assign inp_33[52]=(C[52]|or1) && (R[33]);
  assign inp_33[63:53]=C[63:53] & {11{R[33]&and1}};
  assign inp_34[51:0]=C[51:0] & {52{R[34]}};
  assign inp_34[52]=(C[52]|or1) && (R[34]);
  assign inp_34[63:53]=C[63:53] & {11{R[34]&and1}};
  assign inp_35[51:0]=C[51:0] & {52{R[35]}};
  assign inp_35[52]=(C[52]|or1) && (R[35]);
  assign inp_35[63:53]=C[63:53] & {11{R[35]&and1}};
  assign inp_36[51:0]=C[51:0] & {52{R[36]}};
  assign inp_36[52]=(C[52]|or1) && (R[36]);
  assign inp_36[63:53]=C[63:53] & {11{R[36]&and1}};
  assign inp_37[51:0]=C[51:0] & {52{R[37]}};
  assign inp_37[52]=(C[52]|or1) && (R[37]);
  assign inp_37[63:53]=C[63:53] & {11{R[37]&and1}};
  assign inp_38[51:0]=C[51:0] & {52{R[38]}};
  assign inp_38[52]=(C[52]|or1) && (R[38]);
  assign inp_38[63:53]=C[63:53] & {11{R[38]&and1}};
  assign inp_39[51:0]=C[51:0] & {52{R[39]}};
  assign inp_39[52]=(C[52]|or1) && (R[39]);
  assign inp_39[63:53]=C[63:53] & {11{R[39]&and1}};
  assign inp_40[51:0]=C[51:0] & {52{R[40]}};
  assign inp_40[52]=(C[52]|or1) && (R[40]);
  assign inp_40[63:53]=C[63:53] & {11{R[40]&and1}};
  assign inp_41[51:0]=C[51:0] & {52{R[41]}};
  assign inp_41[52]=(C[52]|or1) && (R[41]);
  assign inp_41[63:53]=C[63:53] & {11{R[41]&and1}};
  assign inp_42[51:0]=C[51:0] & {52{R[42]}};
  assign inp_42[52]=(C[52]|or1) && (R[42]);
  assign inp_42[63:53]=C[63:53] & {11{R[42]&and1}};
  assign inp_43[51:0]=C[51:0] & {52{R[43]}};
  assign inp_43[52]=(C[52]|or1) && (R[43]);
  assign inp_43[63:53]=C[63:53] & {11{R[43]&and1}};
  assign inp_44[51:0]=C[51:0] & {52{R[44]}};
  assign inp_44[52]=(C[52]|or1) && (R[44]);
  assign inp_44[63:53]=C[63:53] & {11{R[44]&and1}};
  assign inp_45[51:0]=C[51:0] & {52{R[45]}};
  assign inp_45[52]=(C[52]|or1) && (R[45]);
  assign inp_45[63:53]=C[63:53] & {11{R[45]&and1}};
  assign inp_46[51:0]=C[51:0] & {52{R[46]}};
  assign inp_46[52]=(C[52]|or1) && (R[46]);
  assign inp_46[63:53]=C[63:53] & {11{R[46]&and1}};
  assign inp_47[51:0]=C[51:0] & {52{R[47]}};
  assign inp_47[52]=(C[52]|or1) && (R[47]);
  assign inp_47[63:53]=C[63:53] & {11{R[47]&and1}};
  assign inp_48[51:0]=C[51:0] & {52{R[48]}};
  assign inp_48[52]=(C[52]|or1) && (R[48]);
  assign inp_48[63:53]=C[63:53] & {11{R[48]&and1}};
  assign inp_49[51:0]=C[51:0] & {52{R[49]}};
  assign inp_49[52]=(C[52]|or1) && (R[49]);
  assign inp_49[63:53]=C[63:53] & {11{R[49]&and1}};
  assign inp_50[51:0]=C[51:0] & {52{R[50]}};
  assign inp_50[52]=(C[52]|or1) && (R[50]);
  assign inp_50[63:53]=C[63:53] & {11{R[50]&and1}};
  assign inp_51[51:0]=C[51:0] & {52{R[51]}};
  assign inp_51[52]=(C[52]|or1) && (R[51]);
  assign inp_51[63:53]=C[63:53] & {11{R[51]&and1}};
  assign inp_52[51:0]=C[51:0] & {52{R[52]|or1}};
  assign inp_52[52]=(C[52]|or1) & (R[52]|or1);
  assign inp_52[63:53]=C[63:53] & {11{R[52]&and1}};
  assign inp_53=C & {64{R[53]&and1}};
  assign inp_54=C & {64{R[54]&and1}};
  assign inp_55=C & {64{R[55]&and1}};
  assign inp_56=C & {64{R[56]&and1}};
  assign inp_57=C & {64{R[57]&and1}};
  assign inp_58=C & {64{R[58]&and1}};
  assign inp_59=C & {64{R[59]&and1}};
  assign inp_60=C & {64{R[60]&and1}};
  assign inp_61=C & {64{R[61]&and1}};
  assign inp_62=C & {64{R[62]&and1}};
  assign inp_63=C & {64{R[63]&and1}};
  assign A_out[0]=REGS_1304;
  assign A_out[1]=REGS_1305;
  assign A_out[2]=REGS_1306;
  assign A_out[3]=REGS_1307;
  assign A_out[4]=REGS_1308;
  assign A_out[5]=REGS_1309;
  assign A_out[6]=REGS_1310;
  assign A_out[7]=REGS_1311;
  assign A_out[8]=REGS_1312;
  assign A_out[9]=HA_out_363;
  assign A_out[10]=HA_out_441;
  assign A_out[11]=HA_cout_441;
  assign A_out[12]=HA_cout_442;
  assign A_out[13]=HA_cout_443;
  assign A_out[14]=HA_cout_444;
  assign A_out[15]=HA_cout_445;
  assign A_out[16]=HA_cout_446;
  assign A_out[17]=HA_cout_447;
  assign A_out[18]=HA_cout_448;
  assign A_out[19]=HA_cout_449;
  assign A_out[20]=HA_cout_450;
  assign A_out[21]=HA_cout_451;
  assign A_out[22]=HA_cout_452;
  assign A_out[23]=HA_cout_453;
  assign A_out[24]=HA_cout_454;
  assign A_out[25]=HA_cout_455;
  assign A_out[26]=HA_cout_456;
  assign A_out[27]=HA_cout_457;
  assign A_out[28]=HA_cout_458;
  assign A_out[29]=HA_cout_459;
  assign A_out[30]=HA_cout_460;
  assign A_out[31]=HA_cout_461;
  assign A_out[32]=HA_cout_462;
  assign A_out[33]=HA_cout_463;
  assign A_out[34]=HA_cout_464;
  assign A_out[35]=HA_cout_465;
  assign A_out[36]=HA_cout_466;
  assign A_out[37]=HA_cout_467;
  assign A_out[38]=HA_cout_468;
  assign A_out[39]=HA_cout_469;
  assign A_out[40]=HA_cout_470;
  assign A_out[41]=HA_cout_471;
  assign A_out[42]=HA_cout_472;
  assign A_out[43]=HA_cout_473;
  assign A_out[44]=HA_cout_474;
  assign A_out[45]=HA_cout_475;
  assign A_out[46]=HA_cout_476;
  assign A_out[47]=HA_cout_477;
  assign A_out[48]=HA_cout_478;
  assign A_out[49]=HA_cout_479;
  assign A_out[50]=HA_cout_480;
  assign A_out[51]=HA_cout_481;
  assign A_out[52]=HA_cout_482;
  assign A_out[53]=HA_cout_483;
  assign A_out[54]=HA_cout_484;
  assign A_out[55]=HA_cout_485;
  assign A_out[56]=HA_cout_486;
  assign A_out[57]=HA_cout_487;
  assign A_out[58]=HA_cout_488;
  assign A_out[59]=HA_cout_489;
  assign A_out[60]=HA_cout_490;
  assign A_out[61]=HA_cout_491;
  assign A_out[62]=HA_cout_492;
  assign A_out[63]=HA_cout_493;
  assign A_out[64]=HA_cout_494;
  assign A_out[65]=HA_cout_495;
  assign A_out[66]=HA_cout_496;
  assign A_out[67]=HA_cout_497;
  assign A_out[68]=FA_cout_3843;
  assign A_out[69]=HA_cout_498;
  assign A_out[70]=HA_cout_499;
  assign A_out[71]=HA_cout_500;
  assign A_out[72]=HA_cout_501;
  assign A_out[73]=HA_cout_502;
  assign B_out[11]=HA_out_442;
  assign B_out[12]=HA_out_443;
  assign B_out[13]=HA_out_444;
  assign B_out[14]=HA_out_445;
  assign B_out[15]=HA_out_446;
  assign B_out[16]=HA_out_447;
  assign B_out[17]=HA_out_448;
  assign B_out[18]=HA_out_449;
  assign B_out[19]=HA_out_450;
  assign B_out[20]=HA_out_451;
  assign B_out[21]=HA_out_452;
  assign B_out[22]=HA_out_453;
  assign B_out[23]=HA_out_454;
  assign B_out[24]=HA_out_455;
  assign B_out[25]=HA_out_456;
  assign B_out[26]=HA_out_457;
  assign B_out[27]=HA_out_458;
  assign B_out[28]=HA_out_459;
  assign B_out[29]=HA_out_460;
  assign B_out[30]=HA_out_461;
  assign B_out[31]=HA_out_462;
  assign B_out[32]=HA_out_463;
  assign B_out[33]=HA_out_464;
  assign B_out[34]=HA_out_465;
  assign B_out[35]=HA_out_466;
  assign B_out[36]=HA_out_467;
  assign B_out[37]=HA_out_468;
  assign B_out[38]=HA_out_469;
  assign B_out[39]=HA_out_470;
  assign B_out[40]=HA_out_471;
  assign B_out[41]=HA_out_472;
  assign B_out[42]=HA_out_473;
  assign B_out[43]=HA_out_474;
  assign B_out[44]=HA_out_475;
  assign B_out[45]=HA_out_476;
  assign B_out[46]=HA_out_477;
  assign B_out[47]=HA_out_478;
  assign B_out[48]=HA_out_479;
  assign B_out[49]=HA_out_480;
  assign B_out[50]=HA_out_481;
  assign B_out[51]=HA_out_482;
  assign B_out[52]=HA_out_483;
  assign B_out[53]=HA_out_484;
  assign B_out[54]=HA_out_485;
  assign B_out[55]=HA_out_486;
  assign B_out[56]=HA_out_487;
  assign B_out[57]=HA_out_488;
  assign B_out[58]=HA_out_489;
  assign B_out[59]=HA_out_490;
  assign B_out[60]=HA_out_491;
  assign B_out[61]=HA_out_492;
  assign B_out[62]=HA_out_493;
  assign B_out[63]=HA_out_494;
  assign B_out[64]=HA_out_495;
  assign B_out[65]=HA_out_496;
  assign B_out[66]=HA_out_497;
  assign B_out[67]=FA_out_3843;
  assign B_out[68]=HA_out_498;
  assign B_out[69]=HA_out_499;
  assign B_out[70]=HA_out_500;
  assign B_out[71]=HA_out_501;
  assign B_out[72]=HA_out_502;
  assign B_out[73]=HA_out_503;
  assign A_out[74]=HA_cout_503;
  assign B_out[74]=HA_out_504;
  assign A_out[75]=HA_cout_504;
  assign B_out[75]=HA_out_505;
  assign A_out[76]=HA_cout_505;
  assign B_out[76]=HA_out_506;
  assign A_out[77]=HA_cout_506;
  assign B_out[77]=HA_out_507;
  assign A_out[78]=HA_cout_507;
  assign B_out[78]=HA_out_508;
  assign A_out[79]=HA_cout_508;
  assign B_out[79]=HA_out_509;
  assign A_out[80]=HA_cout_509;
  assign B_out[80]=HA_out_510;
  assign A_out[81]=HA_cout_510;
  assign B_out[81]=HA_out_511;
  assign A_out[82]=HA_cout_511;
  assign B_out[82]=HA_out_512;
  assign A_out[83]=HA_cout_512;
  assign B_out[83]=HA_out_513;
  assign A_out[84]=HA_cout_513;
  assign B_out[84]=HA_out_514;
  assign A_out[85]=HA_cout_514;
  assign B_out[85]=HA_out_515;
  assign A_out[86]=HA_cout_515;
  assign B_out[86]=HA_out_516;
  assign A_out[87]=HA_cout_516;
  assign B_out[87]=HA_out_517;
  assign A_out[88]=HA_cout_517;
  assign B_out[88]=HA_out_518;
  assign A_out[89]=HA_cout_518;
  assign B_out[89]=HA_out_519;
  assign A_out[90]=HA_cout_519;
  assign B_out[90]=HA_out_520;
  assign A_out[91]=HA_cout_520;
  assign B_out[91]=HA_out_521;
  assign A_out[92]=HA_cout_521;
  assign B_out[92]=HA_out_522;
  assign A_out[93]=HA_cout_522;
  assign B_out[93]=HA_out_523;
  assign A_out[94]=HA_cout_523;
  assign B_out[94]=HA_out_524;
  assign A_out[95]=HA_cout_524;
  assign B_out[95]=HA_out_525;
  assign A_out[96]=HA_cout_525;
  assign B_out[96]=HA_out_526;
  assign A_out[97]=HA_cout_526;
  assign B_out[97]=HA_out_527;
  assign A_out[98]=HA_cout_527;
  assign B_out[98]=HA_out_528;
  assign A_out[99]=HA_cout_528;
  assign B_out[99]=HA_out_529;
  assign A_out[100]=HA_cout_529;
  assign B_out[100]=HA_out_530;
  assign A_out[101]=HA_cout_530;
  assign B_out[101]=HA_out_531;
  assign A_out[102]=HA_cout_531;
  assign B_out[102]=HA_out_532;
  assign A_out[103]=HA_cout_532;
  assign B_out[103]=HA_out_533;
  assign A_out[104]=HA_cout_533;
  assign B_out[104]=HA_out_534;
  assign A_out[105]=HA_cout_534;
  assign B_out[105]=HA_out_535;
  assign A_out[106]=HA_cout_535;
  assign B_out[106]=HA_out_536;
  assign A_out[107]=HA_cout_536;
  assign B_out[107]=HA_out_537;
  assign A_out[108]=HA_cout_537;
  assign B_out[108]=HA_out_538;
  assign A_out[109]=HA_cout_538;
  assign B_out[109]=HA_out_539;
  assign A_out[110]=HA_cout_539;
  assign B_out[110]=HA_out_540;
  assign A_out[111]=HA_cout_540;
  assign B_out[111]=HA_out_541;
  assign A_out[112]=HA_cout_541;
  assign B_out[112]=HA_out_542;
  assign A_out[113]=HA_cout_542;
  assign B_out[113]=HA_out_543;
  assign A_out[114]=HA_cout_543;
  assign B_out[114]=HA_out_544;
  assign A_out[115]=HA_cout_544;
  assign B_out[115]=HA_out_545;
  assign A_out[116]=HA_cout_545;
  assign B_out[116]=HA_out_546;
  assign A_out[117]=HA_cout_546;
  assign B_out[117]=HA_out_547;
  assign A_out[118]=HA_cout_547;
  assign B_out[118]=HA_out_548;
  assign A_out[119]=HA_cout_548;
  assign B_out[119]=HA_out_549;
  assign A_out[120]=HA_cout_549;
  assign B_out[120]=HA_out_550;
  assign A_out[121]=HA_cout_550;
  assign B_out[121]=HA_out_551;
  assign A_out[122]=HA_cout_551;
  assign B_out[122]=HA_out_552;
  assign A_out[123]=HA_cout_552;
  assign B_out[123]=HA_out_553;
  assign A_out[124]=HA_cout_553;
  assign B_out[124]=HA_out_554;
  assign A_out[125]=HA_cout_554;
  assign B_out[125]=HA_out_555;
  assign A_out[126]=HA_cout_555;
  assign B_out[126]=HA_out_556;
  assign A_out[127]=HA_cout_556;
  assign B_out[127]=HA_out_557;
  assign B_out[0]=1'b0;
  assign B_out[1]=1'b0;
  assign B_out[2]=1'b0;
  assign B_out[3]=1'b0;
  assign B_out[4]=1'b0;
  assign B_out[5]=1'b0;
  assign B_out[6]=1'b0;
  assign B_out[7]=1'b0;
  assign B_out[8]=1'b0;
  assign B_out[9]=1'b0;
  assign B_out[10]=1'b0;

  assign {FA_cout_0,FA_out_0}=inp_0[2]+inp_1[1]+inp_2[0];
  assign {FA_cout_1,FA_out_1}=inp_0[3]+inp_1[2]+inp_2[1];
  assign {FA_cout_2,FA_out_2}=inp_0[4]+inp_1[3]+inp_2[2];
  assign {FA_cout_3,FA_out_3}=inp_0[5]+inp_1[4]+inp_2[3];
  assign {FA_cout_4,FA_out_4}=inp_0[6]+inp_1[5]+inp_2[4];
  assign {FA_cout_5,FA_out_5}=inp_0[7]+inp_1[6]+inp_2[5];
  assign {FA_cout_6,FA_out_6}=inp_0[8]+inp_1[7]+inp_2[6];
  assign {FA_cout_7,FA_out_7}=inp_0[9]+inp_1[8]+inp_2[7];
  assign {FA_cout_8,FA_out_8}=inp_0[10]+inp_1[9]+inp_2[8];
  assign {FA_cout_9,FA_out_9}=inp_0[11]+inp_1[10]+inp_2[9];
  assign {FA_cout_10,FA_out_10}=inp_0[12]+inp_1[11]+inp_2[10];
  assign {FA_cout_11,FA_out_11}=inp_0[13]+inp_1[12]+inp_2[11];
  assign {FA_cout_12,FA_out_12}=inp_0[14]+inp_1[13]+inp_2[12];
  assign {FA_cout_13,FA_out_13}=inp_0[15]+inp_1[14]+inp_2[13];
  assign {FA_cout_14,FA_out_14}=inp_0[16]+inp_1[15]+inp_2[14];
  assign {FA_cout_15,FA_out_15}=inp_0[17]+inp_1[16]+inp_2[15];
  assign {FA_cout_16,FA_out_16}=inp_0[18]+inp_1[17]+inp_2[16];
  assign {FA_cout_17,FA_out_17}=inp_0[19]+inp_1[18]+inp_2[17];
  assign {FA_cout_18,FA_out_18}=inp_0[20]+inp_1[19]+inp_2[18];
  assign {FA_cout_19,FA_out_19}=inp_0[21]+inp_1[20]+inp_2[19];
  assign {FA_cout_20,FA_out_20}=inp_0[22]+inp_1[21]+inp_2[20];
  assign {FA_cout_21,FA_out_21}=inp_0[23]+inp_1[22]+inp_2[21];
  assign {FA_cout_22,FA_out_22}=inp_0[24]+inp_1[23]+inp_2[22];
  assign {FA_cout_23,FA_out_23}=inp_0[25]+inp_1[24]+inp_2[23];
  assign {FA_cout_24,FA_out_24}=inp_0[26]+inp_1[25]+inp_2[24];
  assign {FA_cout_25,FA_out_25}=inp_0[27]+inp_1[26]+inp_2[25];
  assign {FA_cout_26,FA_out_26}=inp_0[28]+inp_1[27]+inp_2[26];
  assign {FA_cout_27,FA_out_27}=inp_0[29]+inp_1[28]+inp_2[27];
  assign {FA_cout_28,FA_out_28}=inp_0[30]+inp_1[29]+inp_2[28];
  assign {FA_cout_29,FA_out_29}=inp_0[31]+inp_1[30]+inp_2[29];
  assign {FA_cout_30,FA_out_30}=inp_0[32]+inp_1[31]+inp_2[30];
  assign {FA_cout_31,FA_out_31}=inp_0[33]+inp_1[32]+inp_2[31];
  assign {FA_cout_32,FA_out_32}=inp_0[34]+inp_1[33]+inp_2[32];
  assign {FA_cout_33,FA_out_33}=inp_0[35]+inp_1[34]+inp_2[33];
  assign {FA_cout_34,FA_out_34}=inp_0[36]+inp_1[35]+inp_2[34];
  assign {FA_cout_35,FA_out_35}=inp_0[37]+inp_1[36]+inp_2[35];
  assign {FA_cout_36,FA_out_36}=inp_0[38]+inp_1[37]+inp_2[36];
  assign {FA_cout_37,FA_out_37}=inp_0[39]+inp_1[38]+inp_2[37];
  assign {FA_cout_38,FA_out_38}=inp_0[40]+inp_1[39]+inp_2[38];
  assign {FA_cout_39,FA_out_39}=inp_0[41]+inp_1[40]+inp_2[39];
  assign {FA_cout_40,FA_out_40}=inp_0[42]+inp_1[41]+inp_2[40];
  assign {FA_cout_41,FA_out_41}=inp_0[43]+inp_1[42]+inp_2[41];
  assign {FA_cout_42,FA_out_42}=inp_0[44]+inp_1[43]+inp_2[42];
  assign {FA_cout_43,FA_out_43}=inp_0[45]+inp_1[44]+inp_2[43];
  assign {FA_cout_44,FA_out_44}=inp_0[46]+inp_1[45]+inp_2[44];
  assign {FA_cout_45,FA_out_45}=inp_0[47]+inp_1[46]+inp_2[45];
  assign {FA_cout_46,FA_out_46}=inp_0[48]+inp_1[47]+inp_2[46];
  assign {FA_cout_47,FA_out_47}=inp_0[49]+inp_1[48]+inp_2[47];
  assign {FA_cout_48,FA_out_48}=inp_0[50]+inp_1[49]+inp_2[48];
  assign {FA_cout_49,FA_out_49}=inp_0[51]+inp_1[50]+inp_2[49];
  assign {FA_cout_50,FA_out_50}=inp_0[52]+inp_1[51]+inp_2[50];
  assign {FA_cout_51,FA_out_51}=inp_0[53]+inp_1[52]+inp_2[51];
  assign {FA_cout_52,FA_out_52}=inp_0[54]+inp_1[53]+inp_2[52];
  assign {FA_cout_53,FA_out_53}=inp_0[55]+inp_1[54]+inp_2[53];
  assign {FA_cout_54,FA_out_54}=inp_0[56]+inp_1[55]+inp_2[54];
  assign {FA_cout_55,FA_out_55}=inp_0[57]+inp_1[56]+inp_2[55];
  assign {FA_cout_56,FA_out_56}=inp_0[58]+inp_1[57]+inp_2[56];
  assign {FA_cout_57,FA_out_57}=inp_0[59]+inp_1[58]+inp_2[57];
  assign {FA_cout_58,FA_out_58}=inp_0[60]+inp_1[59]+inp_2[58];
  assign {FA_cout_59,FA_out_59}=inp_0[61]+inp_1[60]+inp_2[59];
  assign {FA_cout_60,FA_out_60}=inp_0[62]+inp_1[61]+inp_2[60];
  assign {FA_cout_61,FA_out_61}=inp_0[63]+inp_1[62]+inp_2[61];
  assign {FA_cout_62,FA_out_62}=inp_1[63]+inp_2[62]+inp_3[61];
  assign {FA_cout_63,FA_out_63}=inp_2[63]+inp_3[62]+inp_4[61];
  assign {FA_cout_64,FA_out_64}=inp_3[2]+inp_4[1]+inp_5[0];
  assign {FA_cout_65,FA_out_65}=inp_3[3]+inp_4[2]+inp_5[1];
  assign {FA_cout_66,FA_out_66}=inp_3[4]+inp_4[3]+inp_5[2];
  assign {FA_cout_67,FA_out_67}=inp_3[5]+inp_4[4]+inp_5[3];
  assign {FA_cout_68,FA_out_68}=inp_3[6]+inp_4[5]+inp_5[4];
  assign {FA_cout_69,FA_out_69}=inp_3[7]+inp_4[6]+inp_5[5];
  assign {FA_cout_70,FA_out_70}=inp_3[8]+inp_4[7]+inp_5[6];
  assign {FA_cout_71,FA_out_71}=inp_3[9]+inp_4[8]+inp_5[7];
  assign {FA_cout_72,FA_out_72}=inp_3[10]+inp_4[9]+inp_5[8];
  assign {FA_cout_73,FA_out_73}=inp_3[11]+inp_4[10]+inp_5[9];
  assign {FA_cout_74,FA_out_74}=inp_3[12]+inp_4[11]+inp_5[10];
  assign {FA_cout_75,FA_out_75}=inp_3[13]+inp_4[12]+inp_5[11];
  assign {FA_cout_76,FA_out_76}=inp_3[14]+inp_4[13]+inp_5[12];
  assign {FA_cout_77,FA_out_77}=inp_3[15]+inp_4[14]+inp_5[13];
  assign {FA_cout_78,FA_out_78}=inp_3[16]+inp_4[15]+inp_5[14];
  assign {FA_cout_79,FA_out_79}=inp_3[17]+inp_4[16]+inp_5[15];
  assign {FA_cout_80,FA_out_80}=inp_3[18]+inp_4[17]+inp_5[16];
  assign {FA_cout_81,FA_out_81}=inp_3[19]+inp_4[18]+inp_5[17];
  assign {FA_cout_82,FA_out_82}=inp_3[20]+inp_4[19]+inp_5[18];
  assign {FA_cout_83,FA_out_83}=inp_3[21]+inp_4[20]+inp_5[19];
  assign {FA_cout_84,FA_out_84}=inp_3[22]+inp_4[21]+inp_5[20];
  assign {FA_cout_85,FA_out_85}=inp_3[23]+inp_4[22]+inp_5[21];
  assign {FA_cout_86,FA_out_86}=inp_3[24]+inp_4[23]+inp_5[22];
  assign {FA_cout_87,FA_out_87}=inp_3[25]+inp_4[24]+inp_5[23];
  assign {FA_cout_88,FA_out_88}=inp_3[26]+inp_4[25]+inp_5[24];
  assign {FA_cout_89,FA_out_89}=inp_3[27]+inp_4[26]+inp_5[25];
  assign {FA_cout_90,FA_out_90}=inp_3[28]+inp_4[27]+inp_5[26];
  assign {FA_cout_91,FA_out_91}=inp_3[29]+inp_4[28]+inp_5[27];
  assign {FA_cout_92,FA_out_92}=inp_3[30]+inp_4[29]+inp_5[28];
  assign {FA_cout_93,FA_out_93}=inp_3[31]+inp_4[30]+inp_5[29];
  assign {FA_cout_94,FA_out_94}=inp_3[32]+inp_4[31]+inp_5[30];
  assign {FA_cout_95,FA_out_95}=inp_3[33]+inp_4[32]+inp_5[31];
  assign {FA_cout_96,FA_out_96}=inp_3[34]+inp_4[33]+inp_5[32];
  assign {FA_cout_97,FA_out_97}=inp_3[35]+inp_4[34]+inp_5[33];
  assign {FA_cout_98,FA_out_98}=inp_3[36]+inp_4[35]+inp_5[34];
  assign {FA_cout_99,FA_out_99}=inp_3[37]+inp_4[36]+inp_5[35];
  assign {FA_cout_100,FA_out_100}=inp_3[38]+inp_4[37]+inp_5[36];
  assign {FA_cout_101,FA_out_101}=inp_3[39]+inp_4[38]+inp_5[37];
  assign {FA_cout_102,FA_out_102}=inp_3[40]+inp_4[39]+inp_5[38];
  assign {FA_cout_103,FA_out_103}=inp_3[41]+inp_4[40]+inp_5[39];
  assign {FA_cout_104,FA_out_104}=inp_3[42]+inp_4[41]+inp_5[40];
  assign {FA_cout_105,FA_out_105}=inp_3[43]+inp_4[42]+inp_5[41];
  assign {FA_cout_106,FA_out_106}=inp_3[44]+inp_4[43]+inp_5[42];
  assign {FA_cout_107,FA_out_107}=inp_3[45]+inp_4[44]+inp_5[43];
  assign {FA_cout_108,FA_out_108}=inp_3[46]+inp_4[45]+inp_5[44];
  assign {FA_cout_109,FA_out_109}=inp_3[47]+inp_4[46]+inp_5[45];
  assign {FA_cout_110,FA_out_110}=inp_3[48]+inp_4[47]+inp_5[46];
  assign {FA_cout_111,FA_out_111}=inp_3[49]+inp_4[48]+inp_5[47];
  assign {FA_cout_112,FA_out_112}=inp_3[50]+inp_4[49]+inp_5[48];
  assign {FA_cout_113,FA_out_113}=inp_3[51]+inp_4[50]+inp_5[49];
  assign {FA_cout_114,FA_out_114}=inp_3[52]+inp_4[51]+inp_5[50];
  assign {FA_cout_115,FA_out_115}=inp_3[53]+inp_4[52]+inp_5[51];
  assign {FA_cout_116,FA_out_116}=inp_3[54]+inp_4[53]+inp_5[52];
  assign {FA_cout_117,FA_out_117}=inp_3[55]+inp_4[54]+inp_5[53];
  assign {FA_cout_118,FA_out_118}=inp_3[56]+inp_4[55]+inp_5[54];
  assign {FA_cout_119,FA_out_119}=inp_3[57]+inp_4[56]+inp_5[55];
  assign {FA_cout_120,FA_out_120}=inp_3[58]+inp_4[57]+inp_5[56];
  assign {FA_cout_121,FA_out_121}=inp_3[59]+inp_4[58]+inp_5[57];
  assign {FA_cout_122,FA_out_122}=inp_3[60]+inp_4[59]+inp_5[58];
  assign {FA_cout_123,FA_out_123}=inp_3[63]+inp_4[62]+inp_5[61];
  assign {FA_cout_124,FA_out_124}=inp_4[60]+inp_5[59]+inp_6[58];
  assign {FA_cout_125,FA_out_125}=inp_4[63]+inp_5[62]+inp_6[61];
  assign {FA_cout_126,FA_out_126}=inp_5[60]+inp_6[59]+inp_7[58];
  assign {FA_cout_127,FA_out_127}=inp_5[63]+inp_6[62]+inp_7[61];
  assign {FA_cout_128,FA_out_128}=inp_6[2]+inp_7[1]+inp_8[0];
  assign {FA_cout_129,FA_out_129}=inp_6[3]+inp_7[2]+inp_8[1];
  assign {FA_cout_130,FA_out_130}=inp_6[4]+inp_7[3]+inp_8[2];
  assign {FA_cout_131,FA_out_131}=inp_6[5]+inp_7[4]+inp_8[3];
  assign {FA_cout_132,FA_out_132}=inp_6[6]+inp_7[5]+inp_8[4];
  assign {FA_cout_133,FA_out_133}=inp_6[7]+inp_7[6]+inp_8[5];
  assign {FA_cout_134,FA_out_134}=inp_6[8]+inp_7[7]+inp_8[6];
  assign {FA_cout_135,FA_out_135}=inp_6[9]+inp_7[8]+inp_8[7];
  assign {FA_cout_136,FA_out_136}=inp_6[10]+inp_7[9]+inp_8[8];
  assign {FA_cout_137,FA_out_137}=inp_6[11]+inp_7[10]+inp_8[9];
  assign {FA_cout_138,FA_out_138}=inp_6[12]+inp_7[11]+inp_8[10];
  assign {FA_cout_139,FA_out_139}=inp_6[13]+inp_7[12]+inp_8[11];
  assign {FA_cout_140,FA_out_140}=inp_6[14]+inp_7[13]+inp_8[12];
  assign {FA_cout_141,FA_out_141}=inp_6[15]+inp_7[14]+inp_8[13];
  assign {FA_cout_142,FA_out_142}=inp_6[16]+inp_7[15]+inp_8[14];
  assign {FA_cout_143,FA_out_143}=inp_6[17]+inp_7[16]+inp_8[15];
  assign {FA_cout_144,FA_out_144}=inp_6[18]+inp_7[17]+inp_8[16];
  assign {FA_cout_145,FA_out_145}=inp_6[19]+inp_7[18]+inp_8[17];
  assign {FA_cout_146,FA_out_146}=inp_6[20]+inp_7[19]+inp_8[18];
  assign {FA_cout_147,FA_out_147}=inp_6[21]+inp_7[20]+inp_8[19];
  assign {FA_cout_148,FA_out_148}=inp_6[22]+inp_7[21]+inp_8[20];
  assign {FA_cout_149,FA_out_149}=inp_6[23]+inp_7[22]+inp_8[21];
  assign {FA_cout_150,FA_out_150}=inp_6[24]+inp_7[23]+inp_8[22];
  assign {FA_cout_151,FA_out_151}=inp_6[25]+inp_7[24]+inp_8[23];
  assign {FA_cout_152,FA_out_152}=inp_6[26]+inp_7[25]+inp_8[24];
  assign {FA_cout_153,FA_out_153}=inp_6[27]+inp_7[26]+inp_8[25];
  assign {FA_cout_154,FA_out_154}=inp_6[28]+inp_7[27]+inp_8[26];
  assign {FA_cout_155,FA_out_155}=inp_6[29]+inp_7[28]+inp_8[27];
  assign {FA_cout_156,FA_out_156}=inp_6[30]+inp_7[29]+inp_8[28];
  assign {FA_cout_157,FA_out_157}=inp_6[31]+inp_7[30]+inp_8[29];
  assign {FA_cout_158,FA_out_158}=inp_6[32]+inp_7[31]+inp_8[30];
  assign {FA_cout_159,FA_out_159}=inp_6[33]+inp_7[32]+inp_8[31];
  assign {FA_cout_160,FA_out_160}=inp_6[34]+inp_7[33]+inp_8[32];
  assign {FA_cout_161,FA_out_161}=inp_6[35]+inp_7[34]+inp_8[33];
  assign {FA_cout_162,FA_out_162}=inp_6[36]+inp_7[35]+inp_8[34];
  assign {FA_cout_163,FA_out_163}=inp_6[37]+inp_7[36]+inp_8[35];
  assign {FA_cout_164,FA_out_164}=inp_6[38]+inp_7[37]+inp_8[36];
  assign {FA_cout_165,FA_out_165}=inp_6[39]+inp_7[38]+inp_8[37];
  assign {FA_cout_166,FA_out_166}=inp_6[40]+inp_7[39]+inp_8[38];
  assign {FA_cout_167,FA_out_167}=inp_6[41]+inp_7[40]+inp_8[39];
  assign {FA_cout_168,FA_out_168}=inp_6[42]+inp_7[41]+inp_8[40];
  assign {FA_cout_169,FA_out_169}=inp_6[43]+inp_7[42]+inp_8[41];
  assign {FA_cout_170,FA_out_170}=inp_6[44]+inp_7[43]+inp_8[42];
  assign {FA_cout_171,FA_out_171}=inp_6[45]+inp_7[44]+inp_8[43];
  assign {FA_cout_172,FA_out_172}=inp_6[46]+inp_7[45]+inp_8[44];
  assign {FA_cout_173,FA_out_173}=inp_6[47]+inp_7[46]+inp_8[45];
  assign {FA_cout_174,FA_out_174}=inp_6[48]+inp_7[47]+inp_8[46];
  assign {FA_cout_175,FA_out_175}=inp_6[49]+inp_7[48]+inp_8[47];
  assign {FA_cout_176,FA_out_176}=inp_6[50]+inp_7[49]+inp_8[48];
  assign {FA_cout_177,FA_out_177}=inp_6[51]+inp_7[50]+inp_8[49];
  assign {FA_cout_178,FA_out_178}=inp_6[52]+inp_7[51]+inp_8[50];
  assign {FA_cout_179,FA_out_179}=inp_6[53]+inp_7[52]+inp_8[51];
  assign {FA_cout_180,FA_out_180}=inp_6[54]+inp_7[53]+inp_8[52];
  assign {FA_cout_181,FA_out_181}=inp_6[55]+inp_7[54]+inp_8[53];
  assign {FA_cout_182,FA_out_182}=inp_6[56]+inp_7[55]+inp_8[54];
  assign {FA_cout_183,FA_out_183}=inp_6[57]+inp_7[56]+inp_8[55];
  assign {FA_cout_184,FA_out_184}=inp_6[60]+inp_7[59]+inp_8[58];
  assign {FA_cout_185,FA_out_185}=inp_6[63]+inp_7[62]+inp_8[61];
  assign {FA_cout_186,FA_out_186}=inp_7[57]+inp_8[56]+inp_9[55];
  assign {FA_cout_187,FA_out_187}=inp_7[60]+inp_8[59]+inp_9[58];
  assign {FA_cout_188,FA_out_188}=inp_7[63]+inp_8[62]+inp_9[61];
  assign {FA_cout_189,FA_out_189}=inp_8[57]+inp_9[56]+inp_10[55];
  assign {FA_cout_190,FA_out_190}=inp_8[60]+inp_9[59]+inp_10[58];
  assign {FA_cout_191,FA_out_191}=inp_8[63]+inp_9[62]+inp_10[61];
  assign {FA_cout_192,FA_out_192}=inp_9[2]+inp_10[1]+inp_11[0];
  assign {FA_cout_193,FA_out_193}=inp_9[3]+inp_10[2]+inp_11[1];
  assign {FA_cout_194,FA_out_194}=inp_9[4]+inp_10[3]+inp_11[2];
  assign {FA_cout_195,FA_out_195}=inp_9[5]+inp_10[4]+inp_11[3];
  assign {FA_cout_196,FA_out_196}=inp_9[6]+inp_10[5]+inp_11[4];
  assign {FA_cout_197,FA_out_197}=inp_9[7]+inp_10[6]+inp_11[5];
  assign {FA_cout_198,FA_out_198}=inp_9[8]+inp_10[7]+inp_11[6];
  assign {FA_cout_199,FA_out_199}=inp_9[9]+inp_10[8]+inp_11[7];
  assign {FA_cout_200,FA_out_200}=inp_9[10]+inp_10[9]+inp_11[8];
  assign {FA_cout_201,FA_out_201}=inp_9[11]+inp_10[10]+inp_11[9];
  assign {FA_cout_202,FA_out_202}=inp_9[12]+inp_10[11]+inp_11[10];
  assign {FA_cout_203,FA_out_203}=inp_9[13]+inp_10[12]+inp_11[11];
  assign {FA_cout_204,FA_out_204}=inp_9[14]+inp_10[13]+inp_11[12];
  assign {FA_cout_205,FA_out_205}=inp_9[15]+inp_10[14]+inp_11[13];
  assign {FA_cout_206,FA_out_206}=inp_9[16]+inp_10[15]+inp_11[14];
  assign {FA_cout_207,FA_out_207}=inp_9[17]+inp_10[16]+inp_11[15];
  assign {FA_cout_208,FA_out_208}=inp_9[18]+inp_10[17]+inp_11[16];
  assign {FA_cout_209,FA_out_209}=inp_9[19]+inp_10[18]+inp_11[17];
  assign {FA_cout_210,FA_out_210}=inp_9[20]+inp_10[19]+inp_11[18];
  assign {FA_cout_211,FA_out_211}=inp_9[21]+inp_10[20]+inp_11[19];
  assign {FA_cout_212,FA_out_212}=inp_9[22]+inp_10[21]+inp_11[20];
  assign {FA_cout_213,FA_out_213}=inp_9[23]+inp_10[22]+inp_11[21];
  assign {FA_cout_214,FA_out_214}=inp_9[24]+inp_10[23]+inp_11[22];
  assign {FA_cout_215,FA_out_215}=inp_9[25]+inp_10[24]+inp_11[23];
  assign {FA_cout_216,FA_out_216}=inp_9[26]+inp_10[25]+inp_11[24];
  assign {FA_cout_217,FA_out_217}=inp_9[27]+inp_10[26]+inp_11[25];
  assign {FA_cout_218,FA_out_218}=inp_9[28]+inp_10[27]+inp_11[26];
  assign {FA_cout_219,FA_out_219}=inp_9[29]+inp_10[28]+inp_11[27];
  assign {FA_cout_220,FA_out_220}=inp_9[30]+inp_10[29]+inp_11[28];
  assign {FA_cout_221,FA_out_221}=inp_9[31]+inp_10[30]+inp_11[29];
  assign {FA_cout_222,FA_out_222}=inp_9[32]+inp_10[31]+inp_11[30];
  assign {FA_cout_223,FA_out_223}=inp_9[33]+inp_10[32]+inp_11[31];
  assign {FA_cout_224,FA_out_224}=inp_9[34]+inp_10[33]+inp_11[32];
  assign {FA_cout_225,FA_out_225}=inp_9[35]+inp_10[34]+inp_11[33];
  assign {FA_cout_226,FA_out_226}=inp_9[36]+inp_10[35]+inp_11[34];
  assign {FA_cout_227,FA_out_227}=inp_9[37]+inp_10[36]+inp_11[35];
  assign {FA_cout_228,FA_out_228}=inp_9[38]+inp_10[37]+inp_11[36];
  assign {FA_cout_229,FA_out_229}=inp_9[39]+inp_10[38]+inp_11[37];
  assign {FA_cout_230,FA_out_230}=inp_9[40]+inp_10[39]+inp_11[38];
  assign {FA_cout_231,FA_out_231}=inp_9[41]+inp_10[40]+inp_11[39];
  assign {FA_cout_232,FA_out_232}=inp_9[42]+inp_10[41]+inp_11[40];
  assign {FA_cout_233,FA_out_233}=inp_9[43]+inp_10[42]+inp_11[41];
  assign {FA_cout_234,FA_out_234}=inp_9[44]+inp_10[43]+inp_11[42];
  assign {FA_cout_235,FA_out_235}=inp_9[45]+inp_10[44]+inp_11[43];
  assign {FA_cout_236,FA_out_236}=inp_9[46]+inp_10[45]+inp_11[44];
  assign {FA_cout_237,FA_out_237}=inp_9[47]+inp_10[46]+inp_11[45];
  assign {FA_cout_238,FA_out_238}=inp_9[48]+inp_10[47]+inp_11[46];
  assign {FA_cout_239,FA_out_239}=inp_9[49]+inp_10[48]+inp_11[47];
  assign {FA_cout_240,FA_out_240}=inp_9[50]+inp_10[49]+inp_11[48];
  assign {FA_cout_241,FA_out_241}=inp_9[51]+inp_10[50]+inp_11[49];
  assign {FA_cout_242,FA_out_242}=inp_9[52]+inp_10[51]+inp_11[50];
  assign {FA_cout_243,FA_out_243}=inp_9[53]+inp_10[52]+inp_11[51];
  assign {FA_cout_244,FA_out_244}=inp_9[54]+inp_10[53]+inp_11[52];
  assign {FA_cout_245,FA_out_245}=inp_9[57]+inp_10[56]+inp_11[55];
  assign {FA_cout_246,FA_out_246}=inp_9[60]+inp_10[59]+inp_11[58];
  assign {FA_cout_247,FA_out_247}=inp_9[63]+inp_10[62]+inp_11[61];
  assign {FA_cout_248,FA_out_248}=inp_10[54]+inp_11[53]+inp_12[52];
  assign {FA_cout_249,FA_out_249}=inp_10[57]+inp_11[56]+inp_12[55];
  assign {FA_cout_250,FA_out_250}=inp_10[60]+inp_11[59]+inp_12[58];
  assign {FA_cout_251,FA_out_251}=inp_10[63]+inp_11[62]+inp_12[61];
  assign {FA_cout_252,FA_out_252}=inp_11[54]+inp_12[53]+inp_13[52];
  assign {FA_cout_253,FA_out_253}=inp_11[57]+inp_12[56]+inp_13[55];
  assign {FA_cout_254,FA_out_254}=inp_11[60]+inp_12[59]+inp_13[58];
  assign {FA_cout_255,FA_out_255}=inp_11[63]+inp_12[62]+inp_13[61];
  assign {FA_cout_256,FA_out_256}=inp_12[2]+inp_13[1]+inp_14[0];
  assign {FA_cout_257,FA_out_257}=inp_12[3]+inp_13[2]+inp_14[1];
  assign {FA_cout_258,FA_out_258}=inp_12[4]+inp_13[3]+inp_14[2];
  assign {FA_cout_259,FA_out_259}=inp_12[5]+inp_13[4]+inp_14[3];
  assign {FA_cout_260,FA_out_260}=inp_12[6]+inp_13[5]+inp_14[4];
  assign {FA_cout_261,FA_out_261}=inp_12[7]+inp_13[6]+inp_14[5];
  assign {FA_cout_262,FA_out_262}=inp_12[8]+inp_13[7]+inp_14[6];
  assign {FA_cout_263,FA_out_263}=inp_12[9]+inp_13[8]+inp_14[7];
  assign {FA_cout_264,FA_out_264}=inp_12[10]+inp_13[9]+inp_14[8];
  assign {FA_cout_265,FA_out_265}=inp_12[11]+inp_13[10]+inp_14[9];
  assign {FA_cout_266,FA_out_266}=inp_12[12]+inp_13[11]+inp_14[10];
  assign {FA_cout_267,FA_out_267}=inp_12[13]+inp_13[12]+inp_14[11];
  assign {FA_cout_268,FA_out_268}=inp_12[14]+inp_13[13]+inp_14[12];
  assign {FA_cout_269,FA_out_269}=inp_12[15]+inp_13[14]+inp_14[13];
  assign {FA_cout_270,FA_out_270}=inp_12[16]+inp_13[15]+inp_14[14];
  assign {FA_cout_271,FA_out_271}=inp_12[17]+inp_13[16]+inp_14[15];
  assign {FA_cout_272,FA_out_272}=inp_12[18]+inp_13[17]+inp_14[16];
  assign {FA_cout_273,FA_out_273}=inp_12[19]+inp_13[18]+inp_14[17];
  assign {FA_cout_274,FA_out_274}=inp_12[20]+inp_13[19]+inp_14[18];
  assign {FA_cout_275,FA_out_275}=inp_12[21]+inp_13[20]+inp_14[19];
  assign {FA_cout_276,FA_out_276}=inp_12[22]+inp_13[21]+inp_14[20];
  assign {FA_cout_277,FA_out_277}=inp_12[23]+inp_13[22]+inp_14[21];
  assign {FA_cout_278,FA_out_278}=inp_12[24]+inp_13[23]+inp_14[22];
  assign {FA_cout_279,FA_out_279}=inp_12[25]+inp_13[24]+inp_14[23];
  assign {FA_cout_280,FA_out_280}=inp_12[26]+inp_13[25]+inp_14[24];
  assign {FA_cout_281,FA_out_281}=inp_12[27]+inp_13[26]+inp_14[25];
  assign {FA_cout_282,FA_out_282}=inp_12[28]+inp_13[27]+inp_14[26];
  assign {FA_cout_283,FA_out_283}=inp_12[29]+inp_13[28]+inp_14[27];
  assign {FA_cout_284,FA_out_284}=inp_12[30]+inp_13[29]+inp_14[28];
  assign {FA_cout_285,FA_out_285}=inp_12[31]+inp_13[30]+inp_14[29];
  assign {FA_cout_286,FA_out_286}=inp_12[32]+inp_13[31]+inp_14[30];
  assign {FA_cout_287,FA_out_287}=inp_12[33]+inp_13[32]+inp_14[31];
  assign {FA_cout_288,FA_out_288}=inp_12[34]+inp_13[33]+inp_14[32];
  assign {FA_cout_289,FA_out_289}=inp_12[35]+inp_13[34]+inp_14[33];
  assign {FA_cout_290,FA_out_290}=inp_12[36]+inp_13[35]+inp_14[34];
  assign {FA_cout_291,FA_out_291}=inp_12[37]+inp_13[36]+inp_14[35];
  assign {FA_cout_292,FA_out_292}=inp_12[38]+inp_13[37]+inp_14[36];
  assign {FA_cout_293,FA_out_293}=inp_12[39]+inp_13[38]+inp_14[37];
  assign {FA_cout_294,FA_out_294}=inp_12[40]+inp_13[39]+inp_14[38];
  assign {FA_cout_295,FA_out_295}=inp_12[41]+inp_13[40]+inp_14[39];
  assign {FA_cout_296,FA_out_296}=inp_12[42]+inp_13[41]+inp_14[40];
  assign {FA_cout_297,FA_out_297}=inp_12[43]+inp_13[42]+inp_14[41];
  assign {FA_cout_298,FA_out_298}=inp_12[44]+inp_13[43]+inp_14[42];
  assign {FA_cout_299,FA_out_299}=inp_12[45]+inp_13[44]+inp_14[43];
  assign {FA_cout_300,FA_out_300}=inp_12[46]+inp_13[45]+inp_14[44];
  assign {FA_cout_301,FA_out_301}=inp_12[47]+inp_13[46]+inp_14[45];
  assign {FA_cout_302,FA_out_302}=inp_12[48]+inp_13[47]+inp_14[46];
  assign {FA_cout_303,FA_out_303}=inp_12[49]+inp_13[48]+inp_14[47];
  assign {FA_cout_304,FA_out_304}=inp_12[50]+inp_13[49]+inp_14[48];
  assign {FA_cout_305,FA_out_305}=inp_12[51]+inp_13[50]+inp_14[49];
  assign {FA_cout_306,FA_out_306}=inp_12[54]+inp_13[53]+inp_14[52];
  assign {FA_cout_307,FA_out_307}=inp_12[57]+inp_13[56]+inp_14[55];
  assign {FA_cout_308,FA_out_308}=inp_12[60]+inp_13[59]+inp_14[58];
  assign {FA_cout_309,FA_out_309}=inp_12[63]+inp_13[62]+inp_14[61];
  assign {FA_cout_310,FA_out_310}=inp_13[51]+inp_14[50]+inp_15[49];
  assign {FA_cout_311,FA_out_311}=inp_13[54]+inp_14[53]+inp_15[52];
  assign {FA_cout_312,FA_out_312}=inp_13[57]+inp_14[56]+inp_15[55];
  assign {FA_cout_313,FA_out_313}=inp_13[60]+inp_14[59]+inp_15[58];
  assign {FA_cout_314,FA_out_314}=inp_13[63]+inp_14[62]+inp_15[61];
  assign {FA_cout_315,FA_out_315}=inp_14[51]+inp_15[50]+inp_16[49];
  assign {FA_cout_316,FA_out_316}=inp_14[54]+inp_15[53]+inp_16[52];
  assign {FA_cout_317,FA_out_317}=inp_14[57]+inp_15[56]+inp_16[55];
  assign {FA_cout_318,FA_out_318}=inp_14[60]+inp_15[59]+inp_16[58];
  assign {FA_cout_319,FA_out_319}=inp_14[63]+inp_15[62]+inp_16[61];
  assign {FA_cout_320,FA_out_320}=inp_15[2]+inp_16[1]+inp_17[0];
  assign {FA_cout_321,FA_out_321}=inp_15[3]+inp_16[2]+inp_17[1];
  assign {FA_cout_322,FA_out_322}=inp_15[4]+inp_16[3]+inp_17[2];
  assign {FA_cout_323,FA_out_323}=inp_15[5]+inp_16[4]+inp_17[3];
  assign {FA_cout_324,FA_out_324}=inp_15[6]+inp_16[5]+inp_17[4];
  assign {FA_cout_325,FA_out_325}=inp_15[7]+inp_16[6]+inp_17[5];
  assign {FA_cout_326,FA_out_326}=inp_15[8]+inp_16[7]+inp_17[6];
  assign {FA_cout_327,FA_out_327}=inp_15[9]+inp_16[8]+inp_17[7];
  assign {FA_cout_328,FA_out_328}=inp_15[10]+inp_16[9]+inp_17[8];
  assign {FA_cout_329,FA_out_329}=inp_15[11]+inp_16[10]+inp_17[9];
  assign {FA_cout_330,FA_out_330}=inp_15[12]+inp_16[11]+inp_17[10];
  assign {FA_cout_331,FA_out_331}=inp_15[13]+inp_16[12]+inp_17[11];
  assign {FA_cout_332,FA_out_332}=inp_15[14]+inp_16[13]+inp_17[12];
  assign {FA_cout_333,FA_out_333}=inp_15[15]+inp_16[14]+inp_17[13];
  assign {FA_cout_334,FA_out_334}=inp_15[16]+inp_16[15]+inp_17[14];
  assign {FA_cout_335,FA_out_335}=inp_15[17]+inp_16[16]+inp_17[15];
  assign {FA_cout_336,FA_out_336}=inp_15[18]+inp_16[17]+inp_17[16];
  assign {FA_cout_337,FA_out_337}=inp_15[19]+inp_16[18]+inp_17[17];
  assign {FA_cout_338,FA_out_338}=inp_15[20]+inp_16[19]+inp_17[18];
  assign {FA_cout_339,FA_out_339}=inp_15[21]+inp_16[20]+inp_17[19];
  assign {FA_cout_340,FA_out_340}=inp_15[22]+inp_16[21]+inp_17[20];
  assign {FA_cout_341,FA_out_341}=inp_15[23]+inp_16[22]+inp_17[21];
  assign {FA_cout_342,FA_out_342}=inp_15[24]+inp_16[23]+inp_17[22];
  assign {FA_cout_343,FA_out_343}=inp_15[25]+inp_16[24]+inp_17[23];
  assign {FA_cout_344,FA_out_344}=inp_15[26]+inp_16[25]+inp_17[24];
  assign {FA_cout_345,FA_out_345}=inp_15[27]+inp_16[26]+inp_17[25];
  assign {FA_cout_346,FA_out_346}=inp_15[28]+inp_16[27]+inp_17[26];
  assign {FA_cout_347,FA_out_347}=inp_15[29]+inp_16[28]+inp_17[27];
  assign {FA_cout_348,FA_out_348}=inp_15[30]+inp_16[29]+inp_17[28];
  assign {FA_cout_349,FA_out_349}=inp_15[31]+inp_16[30]+inp_17[29];
  assign {FA_cout_350,FA_out_350}=inp_15[32]+inp_16[31]+inp_17[30];
  assign {FA_cout_351,FA_out_351}=inp_15[33]+inp_16[32]+inp_17[31];
  assign {FA_cout_352,FA_out_352}=inp_15[34]+inp_16[33]+inp_17[32];
  assign {FA_cout_353,FA_out_353}=inp_15[35]+inp_16[34]+inp_17[33];
  assign {FA_cout_354,FA_out_354}=inp_15[36]+inp_16[35]+inp_17[34];
  assign {FA_cout_355,FA_out_355}=inp_15[37]+inp_16[36]+inp_17[35];
  assign {FA_cout_356,FA_out_356}=inp_15[38]+inp_16[37]+inp_17[36];
  assign {FA_cout_357,FA_out_357}=inp_15[39]+inp_16[38]+inp_17[37];
  assign {FA_cout_358,FA_out_358}=inp_15[40]+inp_16[39]+inp_17[38];
  assign {FA_cout_359,FA_out_359}=inp_15[41]+inp_16[40]+inp_17[39];
  assign {FA_cout_360,FA_out_360}=inp_15[42]+inp_16[41]+inp_17[40];
  assign {FA_cout_361,FA_out_361}=inp_15[43]+inp_16[42]+inp_17[41];
  assign {FA_cout_362,FA_out_362}=inp_15[44]+inp_16[43]+inp_17[42];
  assign {FA_cout_363,FA_out_363}=inp_15[45]+inp_16[44]+inp_17[43];
  assign {FA_cout_364,FA_out_364}=inp_15[46]+inp_16[45]+inp_17[44];
  assign {FA_cout_365,FA_out_365}=inp_15[47]+inp_16[46]+inp_17[45];
  assign {FA_cout_366,FA_out_366}=inp_15[48]+inp_16[47]+inp_17[46];
  assign {FA_cout_367,FA_out_367}=inp_15[51]+inp_16[50]+inp_17[49];
  assign {FA_cout_368,FA_out_368}=inp_15[54]+inp_16[53]+inp_17[52];
  assign {FA_cout_369,FA_out_369}=inp_15[57]+inp_16[56]+inp_17[55];
  assign {FA_cout_370,FA_out_370}=inp_15[60]+inp_16[59]+inp_17[58];
  assign {FA_cout_371,FA_out_371}=inp_15[63]+inp_16[62]+inp_17[61];
  assign {FA_cout_372,FA_out_372}=inp_16[48]+inp_17[47]+inp_18[46];
  assign {FA_cout_373,FA_out_373}=inp_16[51]+inp_17[50]+inp_18[49];
  assign {FA_cout_374,FA_out_374}=inp_16[54]+inp_17[53]+inp_18[52];
  assign {FA_cout_375,FA_out_375}=inp_16[57]+inp_17[56]+inp_18[55];
  assign {FA_cout_376,FA_out_376}=inp_16[60]+inp_17[59]+inp_18[58];
  assign {FA_cout_377,FA_out_377}=inp_16[63]+inp_17[62]+inp_18[61];
  assign {FA_cout_378,FA_out_378}=inp_17[48]+inp_18[47]+inp_19[46];
  assign {FA_cout_379,FA_out_379}=inp_17[51]+inp_18[50]+inp_19[49];
  assign {FA_cout_380,FA_out_380}=inp_17[54]+inp_18[53]+inp_19[52];
  assign {FA_cout_381,FA_out_381}=inp_17[57]+inp_18[56]+inp_19[55];
  assign {FA_cout_382,FA_out_382}=inp_17[60]+inp_18[59]+inp_19[58];
  assign {FA_cout_383,FA_out_383}=inp_17[63]+inp_18[62]+inp_19[61];
  assign {FA_cout_384,FA_out_384}=inp_18[2]+inp_19[1]+inp_20[0];
  assign {FA_cout_385,FA_out_385}=inp_18[3]+inp_19[2]+inp_20[1];
  assign {FA_cout_386,FA_out_386}=inp_18[4]+inp_19[3]+inp_20[2];
  assign {FA_cout_387,FA_out_387}=inp_18[5]+inp_19[4]+inp_20[3];
  assign {FA_cout_388,FA_out_388}=inp_18[6]+inp_19[5]+inp_20[4];
  assign {FA_cout_389,FA_out_389}=inp_18[7]+inp_19[6]+inp_20[5];
  assign {FA_cout_390,FA_out_390}=inp_18[8]+inp_19[7]+inp_20[6];
  assign {FA_cout_391,FA_out_391}=inp_18[9]+inp_19[8]+inp_20[7];
  assign {FA_cout_392,FA_out_392}=inp_18[10]+inp_19[9]+inp_20[8];
  assign {FA_cout_393,FA_out_393}=inp_18[11]+inp_19[10]+inp_20[9];
  assign {FA_cout_394,FA_out_394}=inp_18[12]+inp_19[11]+inp_20[10];
  assign {FA_cout_395,FA_out_395}=inp_18[13]+inp_19[12]+inp_20[11];
  assign {FA_cout_396,FA_out_396}=inp_18[14]+inp_19[13]+inp_20[12];
  assign {FA_cout_397,FA_out_397}=inp_18[15]+inp_19[14]+inp_20[13];
  assign {FA_cout_398,FA_out_398}=inp_18[16]+inp_19[15]+inp_20[14];
  assign {FA_cout_399,FA_out_399}=inp_18[17]+inp_19[16]+inp_20[15];
  assign {FA_cout_400,FA_out_400}=inp_18[18]+inp_19[17]+inp_20[16];
  assign {FA_cout_401,FA_out_401}=inp_18[19]+inp_19[18]+inp_20[17];
  assign {FA_cout_402,FA_out_402}=inp_18[20]+inp_19[19]+inp_20[18];
  assign {FA_cout_403,FA_out_403}=inp_18[21]+inp_19[20]+inp_20[19];
  assign {FA_cout_404,FA_out_404}=inp_18[22]+inp_19[21]+inp_20[20];
  assign {FA_cout_405,FA_out_405}=inp_18[23]+inp_19[22]+inp_20[21];
  assign {FA_cout_406,FA_out_406}=inp_18[24]+inp_19[23]+inp_20[22];
  assign {FA_cout_407,FA_out_407}=inp_18[25]+inp_19[24]+inp_20[23];
  assign {FA_cout_408,FA_out_408}=inp_18[26]+inp_19[25]+inp_20[24];
  assign {FA_cout_409,FA_out_409}=inp_18[27]+inp_19[26]+inp_20[25];
  assign {FA_cout_410,FA_out_410}=inp_18[28]+inp_19[27]+inp_20[26];
  assign {FA_cout_411,FA_out_411}=inp_18[29]+inp_19[28]+inp_20[27];
  assign {FA_cout_412,FA_out_412}=inp_18[30]+inp_19[29]+inp_20[28];
  assign {FA_cout_413,FA_out_413}=inp_18[31]+inp_19[30]+inp_20[29];
  assign {FA_cout_414,FA_out_414}=inp_18[32]+inp_19[31]+inp_20[30];
  assign {FA_cout_415,FA_out_415}=inp_18[33]+inp_19[32]+inp_20[31];
  assign {FA_cout_416,FA_out_416}=inp_18[34]+inp_19[33]+inp_20[32];
  assign {FA_cout_417,FA_out_417}=inp_18[35]+inp_19[34]+inp_20[33];
  assign {FA_cout_418,FA_out_418}=inp_18[36]+inp_19[35]+inp_20[34];
  assign {FA_cout_419,FA_out_419}=inp_18[37]+inp_19[36]+inp_20[35];
  assign {FA_cout_420,FA_out_420}=inp_18[38]+inp_19[37]+inp_20[36];
  assign {FA_cout_421,FA_out_421}=inp_18[39]+inp_19[38]+inp_20[37];
  assign {FA_cout_422,FA_out_422}=inp_18[40]+inp_19[39]+inp_20[38];
  assign {FA_cout_423,FA_out_423}=inp_18[41]+inp_19[40]+inp_20[39];
  assign {FA_cout_424,FA_out_424}=inp_18[42]+inp_19[41]+inp_20[40];
  assign {FA_cout_425,FA_out_425}=inp_18[43]+inp_19[42]+inp_20[41];
  assign {FA_cout_426,FA_out_426}=inp_18[44]+inp_19[43]+inp_20[42];
  assign {FA_cout_427,FA_out_427}=inp_18[45]+inp_19[44]+inp_20[43];
  assign {FA_cout_428,FA_out_428}=inp_18[48]+inp_19[47]+inp_20[46];
  assign {FA_cout_429,FA_out_429}=inp_18[51]+inp_19[50]+inp_20[49];
  assign {FA_cout_430,FA_out_430}=inp_18[54]+inp_19[53]+inp_20[52];
  assign {FA_cout_431,FA_out_431}=inp_18[57]+inp_19[56]+inp_20[55];
  assign {FA_cout_432,FA_out_432}=inp_18[60]+inp_19[59]+inp_20[58];
  assign {FA_cout_433,FA_out_433}=inp_18[63]+inp_19[62]+inp_20[61];
  assign {FA_cout_434,FA_out_434}=inp_19[45]+inp_20[44]+inp_21[43];
  assign {FA_cout_435,FA_out_435}=inp_19[48]+inp_20[47]+inp_21[46];
  assign {FA_cout_436,FA_out_436}=inp_19[51]+inp_20[50]+inp_21[49];
  assign {FA_cout_437,FA_out_437}=inp_19[54]+inp_20[53]+inp_21[52];
  assign {FA_cout_438,FA_out_438}=inp_19[57]+inp_20[56]+inp_21[55];
  assign {FA_cout_439,FA_out_439}=inp_19[60]+inp_20[59]+inp_21[58];
  assign {FA_cout_440,FA_out_440}=inp_19[63]+inp_20[62]+inp_21[61];
  assign {FA_cout_441,FA_out_441}=inp_20[45]+inp_21[44]+inp_22[43];
  assign {FA_cout_442,FA_out_442}=inp_20[48]+inp_21[47]+inp_22[46];
  assign {FA_cout_443,FA_out_443}=inp_20[51]+inp_21[50]+inp_22[49];
  assign {FA_cout_444,FA_out_444}=inp_20[54]+inp_21[53]+inp_22[52];
  assign {FA_cout_445,FA_out_445}=inp_20[57]+inp_21[56]+inp_22[55];
  assign {FA_cout_446,FA_out_446}=inp_20[60]+inp_21[59]+inp_22[58];
  assign {FA_cout_447,FA_out_447}=inp_20[63]+inp_21[62]+inp_22[61];
  assign {FA_cout_448,FA_out_448}=inp_21[2]+inp_22[1]+inp_23[0];
  assign {FA_cout_449,FA_out_449}=inp_21[3]+inp_22[2]+inp_23[1];
  assign {FA_cout_450,FA_out_450}=inp_21[4]+inp_22[3]+inp_23[2];
  assign {FA_cout_451,FA_out_451}=inp_21[5]+inp_22[4]+inp_23[3];
  assign {FA_cout_452,FA_out_452}=inp_21[6]+inp_22[5]+inp_23[4];
  assign {FA_cout_453,FA_out_453}=inp_21[7]+inp_22[6]+inp_23[5];
  assign {FA_cout_454,FA_out_454}=inp_21[8]+inp_22[7]+inp_23[6];
  assign {FA_cout_455,FA_out_455}=inp_21[9]+inp_22[8]+inp_23[7];
  assign {FA_cout_456,FA_out_456}=inp_21[10]+inp_22[9]+inp_23[8];
  assign {FA_cout_457,FA_out_457}=inp_21[11]+inp_22[10]+inp_23[9];
  assign {FA_cout_458,FA_out_458}=inp_21[12]+inp_22[11]+inp_23[10];
  assign {FA_cout_459,FA_out_459}=inp_21[13]+inp_22[12]+inp_23[11];
  assign {FA_cout_460,FA_out_460}=inp_21[14]+inp_22[13]+inp_23[12];
  assign {FA_cout_461,FA_out_461}=inp_21[15]+inp_22[14]+inp_23[13];
  assign {FA_cout_462,FA_out_462}=inp_21[16]+inp_22[15]+inp_23[14];
  assign {FA_cout_463,FA_out_463}=inp_21[17]+inp_22[16]+inp_23[15];
  assign {FA_cout_464,FA_out_464}=inp_21[18]+inp_22[17]+inp_23[16];
  assign {FA_cout_465,FA_out_465}=inp_21[19]+inp_22[18]+inp_23[17];
  assign {FA_cout_466,FA_out_466}=inp_21[20]+inp_22[19]+inp_23[18];
  assign {FA_cout_467,FA_out_467}=inp_21[21]+inp_22[20]+inp_23[19];
  assign {FA_cout_468,FA_out_468}=inp_21[22]+inp_22[21]+inp_23[20];
  assign {FA_cout_469,FA_out_469}=inp_21[23]+inp_22[22]+inp_23[21];
  assign {FA_cout_470,FA_out_470}=inp_21[24]+inp_22[23]+inp_23[22];
  assign {FA_cout_471,FA_out_471}=inp_21[25]+inp_22[24]+inp_23[23];
  assign {FA_cout_472,FA_out_472}=inp_21[26]+inp_22[25]+inp_23[24];
  assign {FA_cout_473,FA_out_473}=inp_21[27]+inp_22[26]+inp_23[25];
  assign {FA_cout_474,FA_out_474}=inp_21[28]+inp_22[27]+inp_23[26];
  assign {FA_cout_475,FA_out_475}=inp_21[29]+inp_22[28]+inp_23[27];
  assign {FA_cout_476,FA_out_476}=inp_21[30]+inp_22[29]+inp_23[28];
  assign {FA_cout_477,FA_out_477}=inp_21[31]+inp_22[30]+inp_23[29];
  assign {FA_cout_478,FA_out_478}=inp_21[32]+inp_22[31]+inp_23[30];
  assign {FA_cout_479,FA_out_479}=inp_21[33]+inp_22[32]+inp_23[31];
  assign {FA_cout_480,FA_out_480}=inp_21[34]+inp_22[33]+inp_23[32];
  assign {FA_cout_481,FA_out_481}=inp_21[35]+inp_22[34]+inp_23[33];
  assign {FA_cout_482,FA_out_482}=inp_21[36]+inp_22[35]+inp_23[34];
  assign {FA_cout_483,FA_out_483}=inp_21[37]+inp_22[36]+inp_23[35];
  assign {FA_cout_484,FA_out_484}=inp_21[38]+inp_22[37]+inp_23[36];
  assign {FA_cout_485,FA_out_485}=inp_21[39]+inp_22[38]+inp_23[37];
  assign {FA_cout_486,FA_out_486}=inp_21[40]+inp_22[39]+inp_23[38];
  assign {FA_cout_487,FA_out_487}=inp_21[41]+inp_22[40]+inp_23[39];
  assign {FA_cout_488,FA_out_488}=inp_21[42]+inp_22[41]+inp_23[40];
  assign {FA_cout_489,FA_out_489}=inp_21[45]+inp_22[44]+inp_23[43];
  assign {FA_cout_490,FA_out_490}=inp_21[48]+inp_22[47]+inp_23[46];
  assign {FA_cout_491,FA_out_491}=inp_21[51]+inp_22[50]+inp_23[49];
  assign {FA_cout_492,FA_out_492}=inp_21[54]+inp_22[53]+inp_23[52];
  assign {FA_cout_493,FA_out_493}=inp_21[57]+inp_22[56]+inp_23[55];
  assign {FA_cout_494,FA_out_494}=inp_21[60]+inp_22[59]+inp_23[58];
  assign {FA_cout_495,FA_out_495}=inp_21[63]+inp_22[62]+inp_23[61];
  assign {FA_cout_496,FA_out_496}=inp_22[42]+inp_23[41]+inp_24[40];
  assign {FA_cout_497,FA_out_497}=inp_22[45]+inp_23[44]+inp_24[43];
  assign {FA_cout_498,FA_out_498}=inp_22[48]+inp_23[47]+inp_24[46];
  assign {FA_cout_499,FA_out_499}=inp_22[51]+inp_23[50]+inp_24[49];
  assign {FA_cout_500,FA_out_500}=inp_22[54]+inp_23[53]+inp_24[52];
  assign {FA_cout_501,FA_out_501}=inp_22[57]+inp_23[56]+inp_24[55];
  assign {FA_cout_502,FA_out_502}=inp_22[60]+inp_23[59]+inp_24[58];
  assign {FA_cout_503,FA_out_503}=inp_22[63]+inp_23[62]+inp_24[61];
  assign {FA_cout_504,FA_out_504}=inp_23[42]+inp_24[41]+inp_25[40];
  assign {FA_cout_505,FA_out_505}=inp_23[45]+inp_24[44]+inp_25[43];
  assign {FA_cout_506,FA_out_506}=inp_23[48]+inp_24[47]+inp_25[46];
  assign {FA_cout_507,FA_out_507}=inp_23[51]+inp_24[50]+inp_25[49];
  assign {FA_cout_508,FA_out_508}=inp_23[54]+inp_24[53]+inp_25[52];
  assign {FA_cout_509,FA_out_509}=inp_23[57]+inp_24[56]+inp_25[55];
  assign {FA_cout_510,FA_out_510}=inp_23[60]+inp_24[59]+inp_25[58];
  assign {FA_cout_511,FA_out_511}=inp_23[63]+inp_24[62]+inp_25[61];
  assign {FA_cout_512,FA_out_512}=inp_24[2]+inp_25[1]+inp_26[0];
  assign {FA_cout_513,FA_out_513}=inp_24[3]+inp_25[2]+inp_26[1];
  assign {FA_cout_514,FA_out_514}=inp_24[4]+inp_25[3]+inp_26[2];
  assign {FA_cout_515,FA_out_515}=inp_24[5]+inp_25[4]+inp_26[3];
  assign {FA_cout_516,FA_out_516}=inp_24[6]+inp_25[5]+inp_26[4];
  assign {FA_cout_517,FA_out_517}=inp_24[7]+inp_25[6]+inp_26[5];
  assign {FA_cout_518,FA_out_518}=inp_24[8]+inp_25[7]+inp_26[6];
  assign {FA_cout_519,FA_out_519}=inp_24[9]+inp_25[8]+inp_26[7];
  assign {FA_cout_520,FA_out_520}=inp_24[10]+inp_25[9]+inp_26[8];
  assign {FA_cout_521,FA_out_521}=inp_24[11]+inp_25[10]+inp_26[9];
  assign {FA_cout_522,FA_out_522}=inp_24[12]+inp_25[11]+inp_26[10];
  assign {FA_cout_523,FA_out_523}=inp_24[13]+inp_25[12]+inp_26[11];
  assign {FA_cout_524,FA_out_524}=inp_24[14]+inp_25[13]+inp_26[12];
  assign {FA_cout_525,FA_out_525}=inp_24[15]+inp_25[14]+inp_26[13];
  assign {FA_cout_526,FA_out_526}=inp_24[16]+inp_25[15]+inp_26[14];
  assign {FA_cout_527,FA_out_527}=inp_24[17]+inp_25[16]+inp_26[15];
  assign {FA_cout_528,FA_out_528}=inp_24[18]+inp_25[17]+inp_26[16];
  assign {FA_cout_529,FA_out_529}=inp_24[19]+inp_25[18]+inp_26[17];
  assign {FA_cout_530,FA_out_530}=inp_24[20]+inp_25[19]+inp_26[18];
  assign {FA_cout_531,FA_out_531}=inp_24[21]+inp_25[20]+inp_26[19];
  assign {FA_cout_532,FA_out_532}=inp_24[22]+inp_25[21]+inp_26[20];
  assign {FA_cout_533,FA_out_533}=inp_24[23]+inp_25[22]+inp_26[21];
  assign {FA_cout_534,FA_out_534}=inp_24[24]+inp_25[23]+inp_26[22];
  assign {FA_cout_535,FA_out_535}=inp_24[25]+inp_25[24]+inp_26[23];
  assign {FA_cout_536,FA_out_536}=inp_24[26]+inp_25[25]+inp_26[24];
  assign {FA_cout_537,FA_out_537}=inp_24[27]+inp_25[26]+inp_26[25];
  assign {FA_cout_538,FA_out_538}=inp_24[28]+inp_25[27]+inp_26[26];
  assign {FA_cout_539,FA_out_539}=inp_24[29]+inp_25[28]+inp_26[27];
  assign {FA_cout_540,FA_out_540}=inp_24[30]+inp_25[29]+inp_26[28];
  assign {FA_cout_541,FA_out_541}=inp_24[31]+inp_25[30]+inp_26[29];
  assign {FA_cout_542,FA_out_542}=inp_24[32]+inp_25[31]+inp_26[30];
  assign {FA_cout_543,FA_out_543}=inp_24[33]+inp_25[32]+inp_26[31];
  assign {FA_cout_544,FA_out_544}=inp_24[34]+inp_25[33]+inp_26[32];
  assign {FA_cout_545,FA_out_545}=inp_24[35]+inp_25[34]+inp_26[33];
  assign {FA_cout_546,FA_out_546}=inp_24[36]+inp_25[35]+inp_26[34];
  assign {FA_cout_547,FA_out_547}=inp_24[37]+inp_25[36]+inp_26[35];
  assign {FA_cout_548,FA_out_548}=inp_24[38]+inp_25[37]+inp_26[36];
  assign {FA_cout_549,FA_out_549}=inp_24[39]+inp_25[38]+inp_26[37];
  assign {FA_cout_550,FA_out_550}=inp_24[42]+inp_25[41]+inp_26[40];
  assign {FA_cout_551,FA_out_551}=inp_24[45]+inp_25[44]+inp_26[43];
  assign {FA_cout_552,FA_out_552}=inp_24[48]+inp_25[47]+inp_26[46];
  assign {FA_cout_553,FA_out_553}=inp_24[51]+inp_25[50]+inp_26[49];
  assign {FA_cout_554,FA_out_554}=inp_24[54]+inp_25[53]+inp_26[52];
  assign {FA_cout_555,FA_out_555}=inp_24[57]+inp_25[56]+inp_26[55];
  assign {FA_cout_556,FA_out_556}=inp_24[60]+inp_25[59]+inp_26[58];
  assign {FA_cout_557,FA_out_557}=inp_24[63]+inp_25[62]+inp_26[61];
  assign {FA_cout_558,FA_out_558}=inp_25[39]+inp_26[38]+inp_27[37];
  assign {FA_cout_559,FA_out_559}=inp_25[42]+inp_26[41]+inp_27[40];
  assign {FA_cout_560,FA_out_560}=inp_25[45]+inp_26[44]+inp_27[43];
  assign {FA_cout_561,FA_out_561}=inp_25[48]+inp_26[47]+inp_27[46];
  assign {FA_cout_562,FA_out_562}=inp_25[51]+inp_26[50]+inp_27[49];
  assign {FA_cout_563,FA_out_563}=inp_25[54]+inp_26[53]+inp_27[52];
  assign {FA_cout_564,FA_out_564}=inp_25[57]+inp_26[56]+inp_27[55];
  assign {FA_cout_565,FA_out_565}=inp_25[60]+inp_26[59]+inp_27[58];
  assign {FA_cout_566,FA_out_566}=inp_25[63]+inp_26[62]+inp_27[61];
  assign {FA_cout_567,FA_out_567}=inp_26[39]+inp_27[38]+inp_28[37];
  assign {FA_cout_568,FA_out_568}=inp_26[42]+inp_27[41]+inp_28[40];
  assign {FA_cout_569,FA_out_569}=inp_26[45]+inp_27[44]+inp_28[43];
  assign {FA_cout_570,FA_out_570}=inp_26[48]+inp_27[47]+inp_28[46];
  assign {FA_cout_571,FA_out_571}=inp_26[51]+inp_27[50]+inp_28[49];
  assign {FA_cout_572,FA_out_572}=inp_26[54]+inp_27[53]+inp_28[52];
  assign {FA_cout_573,FA_out_573}=inp_26[57]+inp_27[56]+inp_28[55];
  assign {FA_cout_574,FA_out_574}=inp_26[60]+inp_27[59]+inp_28[58];
  assign {FA_cout_575,FA_out_575}=inp_26[63]+inp_27[62]+inp_28[61];
  assign {FA_cout_576,FA_out_576}=inp_27[2]+inp_28[1]+inp_29[0];
  assign {FA_cout_577,FA_out_577}=inp_27[3]+inp_28[2]+inp_29[1];
  assign {FA_cout_578,FA_out_578}=inp_27[4]+inp_28[3]+inp_29[2];
  assign {FA_cout_579,FA_out_579}=inp_27[5]+inp_28[4]+inp_29[3];
  assign {FA_cout_580,FA_out_580}=inp_27[6]+inp_28[5]+inp_29[4];
  assign {FA_cout_581,FA_out_581}=inp_27[7]+inp_28[6]+inp_29[5];
  assign {FA_cout_582,FA_out_582}=inp_27[8]+inp_28[7]+inp_29[6];
  assign {FA_cout_583,FA_out_583}=inp_27[9]+inp_28[8]+inp_29[7];
  assign {FA_cout_584,FA_out_584}=inp_27[10]+inp_28[9]+inp_29[8];
  assign {FA_cout_585,FA_out_585}=inp_27[11]+inp_28[10]+inp_29[9];
  assign {FA_cout_586,FA_out_586}=inp_27[12]+inp_28[11]+inp_29[10];
  assign {FA_cout_587,FA_out_587}=inp_27[13]+inp_28[12]+inp_29[11];
  assign {FA_cout_588,FA_out_588}=inp_27[14]+inp_28[13]+inp_29[12];
  assign {FA_cout_589,FA_out_589}=inp_27[15]+inp_28[14]+inp_29[13];
  assign {FA_cout_590,FA_out_590}=inp_27[16]+inp_28[15]+inp_29[14];
  assign {FA_cout_591,FA_out_591}=inp_27[17]+inp_28[16]+inp_29[15];
  assign {FA_cout_592,FA_out_592}=inp_27[18]+inp_28[17]+inp_29[16];
  assign {FA_cout_593,FA_out_593}=inp_27[19]+inp_28[18]+inp_29[17];
  assign {FA_cout_594,FA_out_594}=inp_27[20]+inp_28[19]+inp_29[18];
  assign {FA_cout_595,FA_out_595}=inp_27[21]+inp_28[20]+inp_29[19];
  assign {FA_cout_596,FA_out_596}=inp_27[22]+inp_28[21]+inp_29[20];
  assign {FA_cout_597,FA_out_597}=inp_27[23]+inp_28[22]+inp_29[21];
  assign {FA_cout_598,FA_out_598}=inp_27[24]+inp_28[23]+inp_29[22];
  assign {FA_cout_599,FA_out_599}=inp_27[25]+inp_28[24]+inp_29[23];
  assign {FA_cout_600,FA_out_600}=inp_27[26]+inp_28[25]+inp_29[24];
  assign {FA_cout_601,FA_out_601}=inp_27[27]+inp_28[26]+inp_29[25];
  assign {FA_cout_602,FA_out_602}=inp_27[28]+inp_28[27]+inp_29[26];
  assign {FA_cout_603,FA_out_603}=inp_27[29]+inp_28[28]+inp_29[27];
  assign {FA_cout_604,FA_out_604}=inp_27[30]+inp_28[29]+inp_29[28];
  assign {FA_cout_605,FA_out_605}=inp_27[31]+inp_28[30]+inp_29[29];
  assign {FA_cout_606,FA_out_606}=inp_27[32]+inp_28[31]+inp_29[30];
  assign {FA_cout_607,FA_out_607}=inp_27[33]+inp_28[32]+inp_29[31];
  assign {FA_cout_608,FA_out_608}=inp_27[34]+inp_28[33]+inp_29[32];
  assign {FA_cout_609,FA_out_609}=inp_27[35]+inp_28[34]+inp_29[33];
  assign {FA_cout_610,FA_out_610}=inp_27[36]+inp_28[35]+inp_29[34];
  assign {FA_cout_611,FA_out_611}=inp_27[39]+inp_28[38]+inp_29[37];
  assign {FA_cout_612,FA_out_612}=inp_27[42]+inp_28[41]+inp_29[40];
  assign {FA_cout_613,FA_out_613}=inp_27[45]+inp_28[44]+inp_29[43];
  assign {FA_cout_614,FA_out_614}=inp_27[48]+inp_28[47]+inp_29[46];
  assign {FA_cout_615,FA_out_615}=inp_27[51]+inp_28[50]+inp_29[49];
  assign {FA_cout_616,FA_out_616}=inp_27[54]+inp_28[53]+inp_29[52];
  assign {FA_cout_617,FA_out_617}=inp_27[57]+inp_28[56]+inp_29[55];
  assign {FA_cout_618,FA_out_618}=inp_27[60]+inp_28[59]+inp_29[58];
  assign {FA_cout_619,FA_out_619}=inp_27[63]+inp_28[62]+inp_29[61];
  assign {FA_cout_620,FA_out_620}=inp_28[36]+inp_29[35]+inp_30[34];
  assign {FA_cout_621,FA_out_621}=inp_28[39]+inp_29[38]+inp_30[37];
  assign {FA_cout_622,FA_out_622}=inp_28[42]+inp_29[41]+inp_30[40];
  assign {FA_cout_623,FA_out_623}=inp_28[45]+inp_29[44]+inp_30[43];
  assign {FA_cout_624,FA_out_624}=inp_28[48]+inp_29[47]+inp_30[46];
  assign {FA_cout_625,FA_out_625}=inp_28[51]+inp_29[50]+inp_30[49];
  assign {FA_cout_626,FA_out_626}=inp_28[54]+inp_29[53]+inp_30[52];
  assign {FA_cout_627,FA_out_627}=inp_28[57]+inp_29[56]+inp_30[55];
  assign {FA_cout_628,FA_out_628}=inp_28[60]+inp_29[59]+inp_30[58];
  assign {FA_cout_629,FA_out_629}=inp_28[63]+inp_29[62]+inp_30[61];
  assign {FA_cout_630,FA_out_630}=inp_29[36]+inp_30[35]+inp_31[34];
  assign {FA_cout_631,FA_out_631}=inp_29[39]+inp_30[38]+inp_31[37];
  assign {FA_cout_632,FA_out_632}=inp_29[42]+inp_30[41]+inp_31[40];
  assign {FA_cout_633,FA_out_633}=inp_29[45]+inp_30[44]+inp_31[43];
  assign {FA_cout_634,FA_out_634}=inp_29[48]+inp_30[47]+inp_31[46];
  assign {FA_cout_635,FA_out_635}=inp_29[51]+inp_30[50]+inp_31[49];
  assign {FA_cout_636,FA_out_636}=inp_29[54]+inp_30[53]+inp_31[52];
  assign {FA_cout_637,FA_out_637}=inp_29[57]+inp_30[56]+inp_31[55];
  assign {FA_cout_638,FA_out_638}=inp_29[60]+inp_30[59]+inp_31[58];
  assign {FA_cout_639,FA_out_639}=inp_29[63]+inp_30[62]+inp_31[61];
  assign {FA_cout_640,FA_out_640}=inp_30[2]+inp_31[1]+inp_32[0];
  assign {FA_cout_641,FA_out_641}=inp_30[3]+inp_31[2]+inp_32[1];
  assign {FA_cout_642,FA_out_642}=inp_30[4]+inp_31[3]+inp_32[2];
  assign {FA_cout_643,FA_out_643}=inp_30[5]+inp_31[4]+inp_32[3];
  assign {FA_cout_644,FA_out_644}=inp_30[6]+inp_31[5]+inp_32[4];
  assign {FA_cout_645,FA_out_645}=inp_30[7]+inp_31[6]+inp_32[5];
  assign {FA_cout_646,FA_out_646}=inp_30[8]+inp_31[7]+inp_32[6];
  assign {FA_cout_647,FA_out_647}=inp_30[9]+inp_31[8]+inp_32[7];
  assign {FA_cout_648,FA_out_648}=inp_30[10]+inp_31[9]+inp_32[8];
  assign {FA_cout_649,FA_out_649}=inp_30[11]+inp_31[10]+inp_32[9];
  assign {FA_cout_650,FA_out_650}=inp_30[12]+inp_31[11]+inp_32[10];
  assign {FA_cout_651,FA_out_651}=inp_30[13]+inp_31[12]+inp_32[11];
  assign {FA_cout_652,FA_out_652}=inp_30[14]+inp_31[13]+inp_32[12];
  assign {FA_cout_653,FA_out_653}=inp_30[15]+inp_31[14]+inp_32[13];
  assign {FA_cout_654,FA_out_654}=inp_30[16]+inp_31[15]+inp_32[14];
  assign {FA_cout_655,FA_out_655}=inp_30[17]+inp_31[16]+inp_32[15];
  assign {FA_cout_656,FA_out_656}=inp_30[18]+inp_31[17]+inp_32[16];
  assign {FA_cout_657,FA_out_657}=inp_30[19]+inp_31[18]+inp_32[17];
  assign {FA_cout_658,FA_out_658}=inp_30[20]+inp_31[19]+inp_32[18];
  assign {FA_cout_659,FA_out_659}=inp_30[21]+inp_31[20]+inp_32[19];
  assign {FA_cout_660,FA_out_660}=inp_30[22]+inp_31[21]+inp_32[20];
  assign {FA_cout_661,FA_out_661}=inp_30[23]+inp_31[22]+inp_32[21];
  assign {FA_cout_662,FA_out_662}=inp_30[24]+inp_31[23]+inp_32[22];
  assign {FA_cout_663,FA_out_663}=inp_30[25]+inp_31[24]+inp_32[23];
  assign {FA_cout_664,FA_out_664}=inp_30[26]+inp_31[25]+inp_32[24];
  assign {FA_cout_665,FA_out_665}=inp_30[27]+inp_31[26]+inp_32[25];
  assign {FA_cout_666,FA_out_666}=inp_30[28]+inp_31[27]+inp_32[26];
  assign {FA_cout_667,FA_out_667}=inp_30[29]+inp_31[28]+inp_32[27];
  assign {FA_cout_668,FA_out_668}=inp_30[30]+inp_31[29]+inp_32[28];
  assign {FA_cout_669,FA_out_669}=inp_30[31]+inp_31[30]+inp_32[29];
  assign {FA_cout_670,FA_out_670}=inp_30[32]+inp_31[31]+inp_32[30];
  assign {FA_cout_671,FA_out_671}=inp_30[33]+inp_31[32]+inp_32[31];
  assign {FA_cout_672,FA_out_672}=inp_30[36]+inp_31[35]+inp_32[34];
  assign {FA_cout_673,FA_out_673}=inp_30[39]+inp_31[38]+inp_32[37];
  assign {FA_cout_674,FA_out_674}=inp_30[42]+inp_31[41]+inp_32[40];
  assign {FA_cout_675,FA_out_675}=inp_30[45]+inp_31[44]+inp_32[43];
  assign {FA_cout_676,FA_out_676}=inp_30[48]+inp_31[47]+inp_32[46];
  assign {FA_cout_677,FA_out_677}=inp_30[51]+inp_31[50]+inp_32[49];
  assign {FA_cout_678,FA_out_678}=inp_30[54]+inp_31[53]+inp_32[52];
  assign {FA_cout_679,FA_out_679}=inp_30[57]+inp_31[56]+inp_32[55];
  assign {FA_cout_680,FA_out_680}=inp_30[60]+inp_31[59]+inp_32[58];
  assign {FA_cout_681,FA_out_681}=inp_30[63]+inp_31[62]+inp_32[61];
  assign {FA_cout_682,FA_out_682}=inp_31[33]+inp_32[32]+inp_33[31];
  assign {FA_cout_683,FA_out_683}=inp_31[36]+inp_32[35]+inp_33[34];
  assign {FA_cout_684,FA_out_684}=inp_31[39]+inp_32[38]+inp_33[37];
  assign {FA_cout_685,FA_out_685}=inp_31[42]+inp_32[41]+inp_33[40];
  assign {FA_cout_686,FA_out_686}=inp_31[45]+inp_32[44]+inp_33[43];
  assign {FA_cout_687,FA_out_687}=inp_31[48]+inp_32[47]+inp_33[46];
  assign {FA_cout_688,FA_out_688}=inp_31[51]+inp_32[50]+inp_33[49];
  assign {FA_cout_689,FA_out_689}=inp_31[54]+inp_32[53]+inp_33[52];
  assign {FA_cout_690,FA_out_690}=inp_31[57]+inp_32[56]+inp_33[55];
  assign {FA_cout_691,FA_out_691}=inp_31[60]+inp_32[59]+inp_33[58];
  assign {FA_cout_692,FA_out_692}=inp_31[63]+inp_32[62]+inp_33[61];
  assign {FA_cout_693,FA_out_693}=inp_32[33]+inp_33[32]+inp_34[31];
  assign {FA_cout_694,FA_out_694}=inp_32[36]+inp_33[35]+inp_34[34];
  assign {FA_cout_695,FA_out_695}=inp_32[39]+inp_33[38]+inp_34[37];
  assign {FA_cout_696,FA_out_696}=inp_32[42]+inp_33[41]+inp_34[40];
  assign {FA_cout_697,FA_out_697}=inp_32[45]+inp_33[44]+inp_34[43];
  assign {FA_cout_698,FA_out_698}=inp_32[48]+inp_33[47]+inp_34[46];
  assign {FA_cout_699,FA_out_699}=inp_32[51]+inp_33[50]+inp_34[49];
  assign {FA_cout_700,FA_out_700}=inp_32[54]+inp_33[53]+inp_34[52];
  assign {FA_cout_701,FA_out_701}=inp_32[57]+inp_33[56]+inp_34[55];
  assign {FA_cout_702,FA_out_702}=inp_32[60]+inp_33[59]+inp_34[58];
  assign {FA_cout_703,FA_out_703}=inp_32[63]+inp_33[62]+inp_34[61];
  assign {FA_cout_704,FA_out_704}=inp_33[2]+inp_34[1]+inp_35[0];
  assign {FA_cout_705,FA_out_705}=inp_33[3]+inp_34[2]+inp_35[1];
  assign {FA_cout_706,FA_out_706}=inp_33[4]+inp_34[3]+inp_35[2];
  assign {FA_cout_707,FA_out_707}=inp_33[5]+inp_34[4]+inp_35[3];
  assign {FA_cout_708,FA_out_708}=inp_33[6]+inp_34[5]+inp_35[4];
  assign {FA_cout_709,FA_out_709}=inp_33[7]+inp_34[6]+inp_35[5];
  assign {FA_cout_710,FA_out_710}=inp_33[8]+inp_34[7]+inp_35[6];
  assign {FA_cout_711,FA_out_711}=inp_33[9]+inp_34[8]+inp_35[7];
  assign {FA_cout_712,FA_out_712}=inp_33[10]+inp_34[9]+inp_35[8];
  assign {FA_cout_713,FA_out_713}=inp_33[11]+inp_34[10]+inp_35[9];
  assign {FA_cout_714,FA_out_714}=inp_33[12]+inp_34[11]+inp_35[10];
  assign {FA_cout_715,FA_out_715}=inp_33[13]+inp_34[12]+inp_35[11];
  assign {FA_cout_716,FA_out_716}=inp_33[14]+inp_34[13]+inp_35[12];
  assign {FA_cout_717,FA_out_717}=inp_33[15]+inp_34[14]+inp_35[13];
  assign {FA_cout_718,FA_out_718}=inp_33[16]+inp_34[15]+inp_35[14];
  assign {FA_cout_719,FA_out_719}=inp_33[17]+inp_34[16]+inp_35[15];
  assign {FA_cout_720,FA_out_720}=inp_33[18]+inp_34[17]+inp_35[16];
  assign {FA_cout_721,FA_out_721}=inp_33[19]+inp_34[18]+inp_35[17];
  assign {FA_cout_722,FA_out_722}=inp_33[20]+inp_34[19]+inp_35[18];
  assign {FA_cout_723,FA_out_723}=inp_33[21]+inp_34[20]+inp_35[19];
  assign {FA_cout_724,FA_out_724}=inp_33[22]+inp_34[21]+inp_35[20];
  assign {FA_cout_725,FA_out_725}=inp_33[23]+inp_34[22]+inp_35[21];
  assign {FA_cout_726,FA_out_726}=inp_33[24]+inp_34[23]+inp_35[22];
  assign {FA_cout_727,FA_out_727}=inp_33[25]+inp_34[24]+inp_35[23];
  assign {FA_cout_728,FA_out_728}=inp_33[26]+inp_34[25]+inp_35[24];
  assign {FA_cout_729,FA_out_729}=inp_33[27]+inp_34[26]+inp_35[25];
  assign {FA_cout_730,FA_out_730}=inp_33[28]+inp_34[27]+inp_35[26];
  assign {FA_cout_731,FA_out_731}=inp_33[29]+inp_34[28]+inp_35[27];
  assign {FA_cout_732,FA_out_732}=inp_33[30]+inp_34[29]+inp_35[28];
  assign {FA_cout_733,FA_out_733}=inp_33[33]+inp_34[32]+inp_35[31];
  assign {FA_cout_734,FA_out_734}=inp_33[36]+inp_34[35]+inp_35[34];
  assign {FA_cout_735,FA_out_735}=inp_33[39]+inp_34[38]+inp_35[37];
  assign {FA_cout_736,FA_out_736}=inp_33[42]+inp_34[41]+inp_35[40];
  assign {FA_cout_737,FA_out_737}=inp_33[45]+inp_34[44]+inp_35[43];
  assign {FA_cout_738,FA_out_738}=inp_33[48]+inp_34[47]+inp_35[46];
  assign {FA_cout_739,FA_out_739}=inp_33[51]+inp_34[50]+inp_35[49];
  assign {FA_cout_740,FA_out_740}=inp_33[54]+inp_34[53]+inp_35[52];
  assign {FA_cout_741,FA_out_741}=inp_33[57]+inp_34[56]+inp_35[55];
  assign {FA_cout_742,FA_out_742}=inp_33[60]+inp_34[59]+inp_35[58];
  assign {FA_cout_743,FA_out_743}=inp_33[63]+inp_34[62]+inp_35[61];
  assign {FA_cout_744,FA_out_744}=inp_34[30]+inp_35[29]+inp_36[28];
  assign {FA_cout_745,FA_out_745}=inp_34[33]+inp_35[32]+inp_36[31];
  assign {FA_cout_746,FA_out_746}=inp_34[36]+inp_35[35]+inp_36[34];
  assign {FA_cout_747,FA_out_747}=inp_34[39]+inp_35[38]+inp_36[37];
  assign {FA_cout_748,FA_out_748}=inp_34[42]+inp_35[41]+inp_36[40];
  assign {FA_cout_749,FA_out_749}=inp_34[45]+inp_35[44]+inp_36[43];
  assign {FA_cout_750,FA_out_750}=inp_34[48]+inp_35[47]+inp_36[46];
  assign {FA_cout_751,FA_out_751}=inp_34[51]+inp_35[50]+inp_36[49];
  assign {FA_cout_752,FA_out_752}=inp_34[54]+inp_35[53]+inp_36[52];
  assign {FA_cout_753,FA_out_753}=inp_34[57]+inp_35[56]+inp_36[55];
  assign {FA_cout_754,FA_out_754}=inp_34[60]+inp_35[59]+inp_36[58];
  assign {FA_cout_755,FA_out_755}=inp_34[63]+inp_35[62]+inp_36[61];
  assign {FA_cout_756,FA_out_756}=inp_35[30]+inp_36[29]+inp_37[28];
  assign {FA_cout_757,FA_out_757}=inp_35[33]+inp_36[32]+inp_37[31];
  assign {FA_cout_758,FA_out_758}=inp_35[36]+inp_36[35]+inp_37[34];
  assign {FA_cout_759,FA_out_759}=inp_35[39]+inp_36[38]+inp_37[37];
  assign {FA_cout_760,FA_out_760}=inp_35[42]+inp_36[41]+inp_37[40];
  assign {FA_cout_761,FA_out_761}=inp_35[45]+inp_36[44]+inp_37[43];
  assign {FA_cout_762,FA_out_762}=inp_35[48]+inp_36[47]+inp_37[46];
  assign {FA_cout_763,FA_out_763}=inp_35[51]+inp_36[50]+inp_37[49];
  assign {FA_cout_764,FA_out_764}=inp_35[54]+inp_36[53]+inp_37[52];
  assign {FA_cout_765,FA_out_765}=inp_35[57]+inp_36[56]+inp_37[55];
  assign {FA_cout_766,FA_out_766}=inp_35[60]+inp_36[59]+inp_37[58];
  assign {FA_cout_767,FA_out_767}=inp_35[63]+inp_36[62]+inp_37[61];
  assign {FA_cout_768,FA_out_768}=inp_36[2]+inp_37[1]+inp_38[0];
  assign {FA_cout_769,FA_out_769}=inp_36[3]+inp_37[2]+inp_38[1];
  assign {FA_cout_770,FA_out_770}=inp_36[4]+inp_37[3]+inp_38[2];
  assign {FA_cout_771,FA_out_771}=inp_36[5]+inp_37[4]+inp_38[3];
  assign {FA_cout_772,FA_out_772}=inp_36[6]+inp_37[5]+inp_38[4];
  assign {FA_cout_773,FA_out_773}=inp_36[7]+inp_37[6]+inp_38[5];
  assign {FA_cout_774,FA_out_774}=inp_36[8]+inp_37[7]+inp_38[6];
  assign {FA_cout_775,FA_out_775}=inp_36[9]+inp_37[8]+inp_38[7];
  assign {FA_cout_776,FA_out_776}=inp_36[10]+inp_37[9]+inp_38[8];
  assign {FA_cout_777,FA_out_777}=inp_36[11]+inp_37[10]+inp_38[9];
  assign {FA_cout_778,FA_out_778}=inp_36[12]+inp_37[11]+inp_38[10];
  assign {FA_cout_779,FA_out_779}=inp_36[13]+inp_37[12]+inp_38[11];
  assign {FA_cout_780,FA_out_780}=inp_36[14]+inp_37[13]+inp_38[12];
  assign {FA_cout_781,FA_out_781}=inp_36[15]+inp_37[14]+inp_38[13];
  assign {FA_cout_782,FA_out_782}=inp_36[16]+inp_37[15]+inp_38[14];
  assign {FA_cout_783,FA_out_783}=inp_36[17]+inp_37[16]+inp_38[15];
  assign {FA_cout_784,FA_out_784}=inp_36[18]+inp_37[17]+inp_38[16];
  assign {FA_cout_785,FA_out_785}=inp_36[19]+inp_37[18]+inp_38[17];
  assign {FA_cout_786,FA_out_786}=inp_36[20]+inp_37[19]+inp_38[18];
  assign {FA_cout_787,FA_out_787}=inp_36[21]+inp_37[20]+inp_38[19];
  assign {FA_cout_788,FA_out_788}=inp_36[22]+inp_37[21]+inp_38[20];
  assign {FA_cout_789,FA_out_789}=inp_36[23]+inp_37[22]+inp_38[21];
  assign {FA_cout_790,FA_out_790}=inp_36[24]+inp_37[23]+inp_38[22];
  assign {FA_cout_791,FA_out_791}=inp_36[25]+inp_37[24]+inp_38[23];
  assign {FA_cout_792,FA_out_792}=inp_36[26]+inp_37[25]+inp_38[24];
  assign {FA_cout_793,FA_out_793}=inp_36[27]+inp_37[26]+inp_38[25];
  assign {FA_cout_794,FA_out_794}=inp_36[30]+inp_37[29]+inp_38[28];
  assign {FA_cout_795,FA_out_795}=inp_36[33]+inp_37[32]+inp_38[31];
  assign {FA_cout_796,FA_out_796}=inp_36[36]+inp_37[35]+inp_38[34];
  assign {FA_cout_797,FA_out_797}=inp_36[39]+inp_37[38]+inp_38[37];
  assign {FA_cout_798,FA_out_798}=inp_36[42]+inp_37[41]+inp_38[40];
  assign {FA_cout_799,FA_out_799}=inp_36[45]+inp_37[44]+inp_38[43];
  assign {FA_cout_800,FA_out_800}=inp_36[48]+inp_37[47]+inp_38[46];
  assign {FA_cout_801,FA_out_801}=inp_36[51]+inp_37[50]+inp_38[49];
  assign {FA_cout_802,FA_out_802}=inp_36[54]+inp_37[53]+inp_38[52];
  assign {FA_cout_803,FA_out_803}=inp_36[57]+inp_37[56]+inp_38[55];
  assign {FA_cout_804,FA_out_804}=inp_36[60]+inp_37[59]+inp_38[58];
  assign {FA_cout_805,FA_out_805}=inp_36[63]+inp_37[62]+inp_38[61];
  assign {FA_cout_806,FA_out_806}=inp_37[27]+inp_38[26]+inp_39[25];
  assign {FA_cout_807,FA_out_807}=inp_37[30]+inp_38[29]+inp_39[28];
  assign {FA_cout_808,FA_out_808}=inp_37[33]+inp_38[32]+inp_39[31];
  assign {FA_cout_809,FA_out_809}=inp_37[36]+inp_38[35]+inp_39[34];
  assign {FA_cout_810,FA_out_810}=inp_37[39]+inp_38[38]+inp_39[37];
  assign {FA_cout_811,FA_out_811}=inp_37[42]+inp_38[41]+inp_39[40];
  assign {FA_cout_812,FA_out_812}=inp_37[45]+inp_38[44]+inp_39[43];
  assign {FA_cout_813,FA_out_813}=inp_37[48]+inp_38[47]+inp_39[46];
  assign {FA_cout_814,FA_out_814}=inp_37[51]+inp_38[50]+inp_39[49];
  assign {FA_cout_815,FA_out_815}=inp_37[54]+inp_38[53]+inp_39[52];
  assign {FA_cout_816,FA_out_816}=inp_37[57]+inp_38[56]+inp_39[55];
  assign {FA_cout_817,FA_out_817}=inp_37[60]+inp_38[59]+inp_39[58];
  assign {FA_cout_818,FA_out_818}=inp_37[63]+inp_38[62]+inp_39[61];
  assign {FA_cout_819,FA_out_819}=inp_38[27]+inp_39[26]+inp_40[25];
  assign {FA_cout_820,FA_out_820}=inp_38[30]+inp_39[29]+inp_40[28];
  assign {FA_cout_821,FA_out_821}=inp_38[33]+inp_39[32]+inp_40[31];
  assign {FA_cout_822,FA_out_822}=inp_38[36]+inp_39[35]+inp_40[34];
  assign {FA_cout_823,FA_out_823}=inp_38[39]+inp_39[38]+inp_40[37];
  assign {FA_cout_824,FA_out_824}=inp_38[42]+inp_39[41]+inp_40[40];
  assign {FA_cout_825,FA_out_825}=inp_38[45]+inp_39[44]+inp_40[43];
  assign {FA_cout_826,FA_out_826}=inp_38[48]+inp_39[47]+inp_40[46];
  assign {FA_cout_827,FA_out_827}=inp_38[51]+inp_39[50]+inp_40[49];
  assign {FA_cout_828,FA_out_828}=inp_38[54]+inp_39[53]+inp_40[52];
  assign {FA_cout_829,FA_out_829}=inp_38[57]+inp_39[56]+inp_40[55];
  assign {FA_cout_830,FA_out_830}=inp_38[60]+inp_39[59]+inp_40[58];
  assign {FA_cout_831,FA_out_831}=inp_38[63]+inp_39[62]+inp_40[61];
  assign {FA_cout_832,FA_out_832}=inp_39[2]+inp_40[1]+inp_41[0];
  assign {FA_cout_833,FA_out_833}=inp_39[3]+inp_40[2]+inp_41[1];
  assign {FA_cout_834,FA_out_834}=inp_39[4]+inp_40[3]+inp_41[2];
  assign {FA_cout_835,FA_out_835}=inp_39[5]+inp_40[4]+inp_41[3];
  assign {FA_cout_836,FA_out_836}=inp_39[6]+inp_40[5]+inp_41[4];
  assign {FA_cout_837,FA_out_837}=inp_39[7]+inp_40[6]+inp_41[5];
  assign {FA_cout_838,FA_out_838}=inp_39[8]+inp_40[7]+inp_41[6];
  assign {FA_cout_839,FA_out_839}=inp_39[9]+inp_40[8]+inp_41[7];
  assign {FA_cout_840,FA_out_840}=inp_39[10]+inp_40[9]+inp_41[8];
  assign {FA_cout_841,FA_out_841}=inp_39[11]+inp_40[10]+inp_41[9];
  assign {FA_cout_842,FA_out_842}=inp_39[12]+inp_40[11]+inp_41[10];
  assign {FA_cout_843,FA_out_843}=inp_39[13]+inp_40[12]+inp_41[11];
  assign {FA_cout_844,FA_out_844}=inp_39[14]+inp_40[13]+inp_41[12];
  assign {FA_cout_845,FA_out_845}=inp_39[15]+inp_40[14]+inp_41[13];
  assign {FA_cout_846,FA_out_846}=inp_39[16]+inp_40[15]+inp_41[14];
  assign {FA_cout_847,FA_out_847}=inp_39[17]+inp_40[16]+inp_41[15];
  assign {FA_cout_848,FA_out_848}=inp_39[18]+inp_40[17]+inp_41[16];
  assign {FA_cout_849,FA_out_849}=inp_39[19]+inp_40[18]+inp_41[17];
  assign {FA_cout_850,FA_out_850}=inp_39[20]+inp_40[19]+inp_41[18];
  assign {FA_cout_851,FA_out_851}=inp_39[21]+inp_40[20]+inp_41[19];
  assign {FA_cout_852,FA_out_852}=inp_39[22]+inp_40[21]+inp_41[20];
  assign {FA_cout_853,FA_out_853}=inp_39[23]+inp_40[22]+inp_41[21];
  assign {FA_cout_854,FA_out_854}=inp_39[24]+inp_40[23]+inp_41[22];
  assign {FA_cout_855,FA_out_855}=inp_39[27]+inp_40[26]+inp_41[25];
  assign {FA_cout_856,FA_out_856}=inp_39[30]+inp_40[29]+inp_41[28];
  assign {FA_cout_857,FA_out_857}=inp_39[33]+inp_40[32]+inp_41[31];
  assign {FA_cout_858,FA_out_858}=inp_39[36]+inp_40[35]+inp_41[34];
  assign {FA_cout_859,FA_out_859}=inp_39[39]+inp_40[38]+inp_41[37];
  assign {FA_cout_860,FA_out_860}=inp_39[42]+inp_40[41]+inp_41[40];
  assign {FA_cout_861,FA_out_861}=inp_39[45]+inp_40[44]+inp_41[43];
  assign {FA_cout_862,FA_out_862}=inp_39[48]+inp_40[47]+inp_41[46];
  assign {FA_cout_863,FA_out_863}=inp_39[51]+inp_40[50]+inp_41[49];
  assign {FA_cout_864,FA_out_864}=inp_39[54]+inp_40[53]+inp_41[52];
  assign {FA_cout_865,FA_out_865}=inp_39[57]+inp_40[56]+inp_41[55];
  assign {FA_cout_866,FA_out_866}=inp_39[60]+inp_40[59]+inp_41[58];
  assign {FA_cout_867,FA_out_867}=inp_39[63]+inp_40[62]+inp_41[61];
  assign {FA_cout_868,FA_out_868}=inp_40[24]+inp_41[23]+inp_42[22];
  assign {FA_cout_869,FA_out_869}=inp_40[27]+inp_41[26]+inp_42[25];
  assign {FA_cout_870,FA_out_870}=inp_40[30]+inp_41[29]+inp_42[28];
  assign {FA_cout_871,FA_out_871}=inp_40[33]+inp_41[32]+inp_42[31];
  assign {FA_cout_872,FA_out_872}=inp_40[36]+inp_41[35]+inp_42[34];
  assign {FA_cout_873,FA_out_873}=inp_40[39]+inp_41[38]+inp_42[37];
  assign {FA_cout_874,FA_out_874}=inp_40[42]+inp_41[41]+inp_42[40];
  assign {FA_cout_875,FA_out_875}=inp_40[45]+inp_41[44]+inp_42[43];
  assign {FA_cout_876,FA_out_876}=inp_40[48]+inp_41[47]+inp_42[46];
  assign {FA_cout_877,FA_out_877}=inp_40[51]+inp_41[50]+inp_42[49];
  assign {FA_cout_878,FA_out_878}=inp_40[54]+inp_41[53]+inp_42[52];
  assign {FA_cout_879,FA_out_879}=inp_40[57]+inp_41[56]+inp_42[55];
  assign {FA_cout_880,FA_out_880}=inp_40[60]+inp_41[59]+inp_42[58];
  assign {FA_cout_881,FA_out_881}=inp_40[63]+inp_41[62]+inp_42[61];
  assign {FA_cout_882,FA_out_882}=inp_41[24]+inp_42[23]+inp_43[22];
  assign {FA_cout_883,FA_out_883}=inp_41[27]+inp_42[26]+inp_43[25];
  assign {FA_cout_884,FA_out_884}=inp_41[30]+inp_42[29]+inp_43[28];
  assign {FA_cout_885,FA_out_885}=inp_41[33]+inp_42[32]+inp_43[31];
  assign {FA_cout_886,FA_out_886}=inp_41[36]+inp_42[35]+inp_43[34];
  assign {FA_cout_887,FA_out_887}=inp_41[39]+inp_42[38]+inp_43[37];
  assign {FA_cout_888,FA_out_888}=inp_41[42]+inp_42[41]+inp_43[40];
  assign {FA_cout_889,FA_out_889}=inp_41[45]+inp_42[44]+inp_43[43];
  assign {FA_cout_890,FA_out_890}=inp_41[48]+inp_42[47]+inp_43[46];
  assign {FA_cout_891,FA_out_891}=inp_41[51]+inp_42[50]+inp_43[49];
  assign {FA_cout_892,FA_out_892}=inp_41[54]+inp_42[53]+inp_43[52];
  assign {FA_cout_893,FA_out_893}=inp_41[57]+inp_42[56]+inp_43[55];
  assign {FA_cout_894,FA_out_894}=inp_41[60]+inp_42[59]+inp_43[58];
  assign {FA_cout_895,FA_out_895}=inp_41[63]+inp_42[62]+inp_43[61];
  assign {FA_cout_896,FA_out_896}=inp_42[2]+inp_43[1]+inp_44[0];
  assign {FA_cout_897,FA_out_897}=inp_42[3]+inp_43[2]+inp_44[1];
  assign {FA_cout_898,FA_out_898}=inp_42[4]+inp_43[3]+inp_44[2];
  assign {FA_cout_899,FA_out_899}=inp_42[5]+inp_43[4]+inp_44[3];
  assign {FA_cout_900,FA_out_900}=inp_42[6]+inp_43[5]+inp_44[4];
  assign {FA_cout_901,FA_out_901}=inp_42[7]+inp_43[6]+inp_44[5];
  assign {FA_cout_902,FA_out_902}=inp_42[8]+inp_43[7]+inp_44[6];
  assign {FA_cout_903,FA_out_903}=inp_42[9]+inp_43[8]+inp_44[7];
  assign {FA_cout_904,FA_out_904}=inp_42[10]+inp_43[9]+inp_44[8];
  assign {FA_cout_905,FA_out_905}=inp_42[11]+inp_43[10]+inp_44[9];
  assign {FA_cout_906,FA_out_906}=inp_42[12]+inp_43[11]+inp_44[10];
  assign {FA_cout_907,FA_out_907}=inp_42[13]+inp_43[12]+inp_44[11];
  assign {FA_cout_908,FA_out_908}=inp_42[14]+inp_43[13]+inp_44[12];
  assign {FA_cout_909,FA_out_909}=inp_42[15]+inp_43[14]+inp_44[13];
  assign {FA_cout_910,FA_out_910}=inp_42[16]+inp_43[15]+inp_44[14];
  assign {FA_cout_911,FA_out_911}=inp_42[17]+inp_43[16]+inp_44[15];
  assign {FA_cout_912,FA_out_912}=inp_42[18]+inp_43[17]+inp_44[16];
  assign {FA_cout_913,FA_out_913}=inp_42[19]+inp_43[18]+inp_44[17];
  assign {FA_cout_914,FA_out_914}=inp_42[20]+inp_43[19]+inp_44[18];
  assign {FA_cout_915,FA_out_915}=inp_42[21]+inp_43[20]+inp_44[19];
  assign {FA_cout_916,FA_out_916}=inp_42[24]+inp_43[23]+inp_44[22];
  assign {FA_cout_917,FA_out_917}=inp_42[27]+inp_43[26]+inp_44[25];
  assign {FA_cout_918,FA_out_918}=inp_42[30]+inp_43[29]+inp_44[28];
  assign {FA_cout_919,FA_out_919}=inp_42[33]+inp_43[32]+inp_44[31];
  assign {FA_cout_920,FA_out_920}=inp_42[36]+inp_43[35]+inp_44[34];
  assign {FA_cout_921,FA_out_921}=inp_42[39]+inp_43[38]+inp_44[37];
  assign {FA_cout_922,FA_out_922}=inp_42[42]+inp_43[41]+inp_44[40];
  assign {FA_cout_923,FA_out_923}=inp_42[45]+inp_43[44]+inp_44[43];
  assign {FA_cout_924,FA_out_924}=inp_42[48]+inp_43[47]+inp_44[46];
  assign {FA_cout_925,FA_out_925}=inp_42[51]+inp_43[50]+inp_44[49];
  assign {FA_cout_926,FA_out_926}=inp_42[54]+inp_43[53]+inp_44[52];
  assign {FA_cout_927,FA_out_927}=inp_42[57]+inp_43[56]+inp_44[55];
  assign {FA_cout_928,FA_out_928}=inp_42[60]+inp_43[59]+inp_44[58];
  assign {FA_cout_929,FA_out_929}=inp_42[63]+inp_43[62]+inp_44[61];
  assign {FA_cout_930,FA_out_930}=inp_43[21]+inp_44[20]+inp_45[19];
  assign {FA_cout_931,FA_out_931}=inp_43[24]+inp_44[23]+inp_45[22];
  assign {FA_cout_932,FA_out_932}=inp_43[27]+inp_44[26]+inp_45[25];
  assign {FA_cout_933,FA_out_933}=inp_43[30]+inp_44[29]+inp_45[28];
  assign {FA_cout_934,FA_out_934}=inp_43[33]+inp_44[32]+inp_45[31];
  assign {FA_cout_935,FA_out_935}=inp_43[36]+inp_44[35]+inp_45[34];
  assign {FA_cout_936,FA_out_936}=inp_43[39]+inp_44[38]+inp_45[37];
  assign {FA_cout_937,FA_out_937}=inp_43[42]+inp_44[41]+inp_45[40];
  assign {FA_cout_938,FA_out_938}=inp_43[45]+inp_44[44]+inp_45[43];
  assign {FA_cout_939,FA_out_939}=inp_43[48]+inp_44[47]+inp_45[46];
  assign {FA_cout_940,FA_out_940}=inp_43[51]+inp_44[50]+inp_45[49];
  assign {FA_cout_941,FA_out_941}=inp_43[54]+inp_44[53]+inp_45[52];
  assign {FA_cout_942,FA_out_942}=inp_43[57]+inp_44[56]+inp_45[55];
  assign {FA_cout_943,FA_out_943}=inp_43[60]+inp_44[59]+inp_45[58];
  assign {FA_cout_944,FA_out_944}=inp_43[63]+inp_44[62]+inp_45[61];
  assign {FA_cout_945,FA_out_945}=inp_44[21]+inp_45[20]+inp_46[19];
  assign {FA_cout_946,FA_out_946}=inp_44[24]+inp_45[23]+inp_46[22];
  assign {FA_cout_947,FA_out_947}=inp_44[27]+inp_45[26]+inp_46[25];
  assign {FA_cout_948,FA_out_948}=inp_44[30]+inp_45[29]+inp_46[28];
  assign {FA_cout_949,FA_out_949}=inp_44[33]+inp_45[32]+inp_46[31];
  assign {FA_cout_950,FA_out_950}=inp_44[36]+inp_45[35]+inp_46[34];
  assign {FA_cout_951,FA_out_951}=inp_44[39]+inp_45[38]+inp_46[37];
  assign {FA_cout_952,FA_out_952}=inp_44[42]+inp_45[41]+inp_46[40];
  assign {FA_cout_953,FA_out_953}=inp_44[45]+inp_45[44]+inp_46[43];
  assign {FA_cout_954,FA_out_954}=inp_44[48]+inp_45[47]+inp_46[46];
  assign {FA_cout_955,FA_out_955}=inp_44[51]+inp_45[50]+inp_46[49];
  assign {FA_cout_956,FA_out_956}=inp_44[54]+inp_45[53]+inp_46[52];
  assign {FA_cout_957,FA_out_957}=inp_44[57]+inp_45[56]+inp_46[55];
  assign {FA_cout_958,FA_out_958}=inp_44[60]+inp_45[59]+inp_46[58];
  assign {FA_cout_959,FA_out_959}=inp_44[63]+inp_45[62]+inp_46[61];
  assign {FA_cout_960,FA_out_960}=inp_45[2]+inp_46[1]+inp_47[0];
  assign {FA_cout_961,FA_out_961}=inp_45[3]+inp_46[2]+inp_47[1];
  assign {FA_cout_962,FA_out_962}=inp_45[4]+inp_46[3]+inp_47[2];
  assign {FA_cout_963,FA_out_963}=inp_45[5]+inp_46[4]+inp_47[3];
  assign {FA_cout_964,FA_out_964}=inp_45[6]+inp_46[5]+inp_47[4];
  assign {FA_cout_965,FA_out_965}=inp_45[7]+inp_46[6]+inp_47[5];
  assign {FA_cout_966,FA_out_966}=inp_45[8]+inp_46[7]+inp_47[6];
  assign {FA_cout_967,FA_out_967}=inp_45[9]+inp_46[8]+inp_47[7];
  assign {FA_cout_968,FA_out_968}=inp_45[10]+inp_46[9]+inp_47[8];
  assign {FA_cout_969,FA_out_969}=inp_45[11]+inp_46[10]+inp_47[9];
  assign {FA_cout_970,FA_out_970}=inp_45[12]+inp_46[11]+inp_47[10];
  assign {FA_cout_971,FA_out_971}=inp_45[13]+inp_46[12]+inp_47[11];
  assign {FA_cout_972,FA_out_972}=inp_45[14]+inp_46[13]+inp_47[12];
  assign {FA_cout_973,FA_out_973}=inp_45[15]+inp_46[14]+inp_47[13];
  assign {FA_cout_974,FA_out_974}=inp_45[16]+inp_46[15]+inp_47[14];
  assign {FA_cout_975,FA_out_975}=inp_45[17]+inp_46[16]+inp_47[15];
  assign {FA_cout_976,FA_out_976}=inp_45[18]+inp_46[17]+inp_47[16];
  assign {FA_cout_977,FA_out_977}=inp_45[21]+inp_46[20]+inp_47[19];
  assign {FA_cout_978,FA_out_978}=inp_45[24]+inp_46[23]+inp_47[22];
  assign {FA_cout_979,FA_out_979}=inp_45[27]+inp_46[26]+inp_47[25];
  assign {FA_cout_980,FA_out_980}=inp_45[30]+inp_46[29]+inp_47[28];
  assign {FA_cout_981,FA_out_981}=inp_45[33]+inp_46[32]+inp_47[31];
  assign {FA_cout_982,FA_out_982}=inp_45[36]+inp_46[35]+inp_47[34];
  assign {FA_cout_983,FA_out_983}=inp_45[39]+inp_46[38]+inp_47[37];
  assign {FA_cout_984,FA_out_984}=inp_45[42]+inp_46[41]+inp_47[40];
  assign {FA_cout_985,FA_out_985}=inp_45[45]+inp_46[44]+inp_47[43];
  assign {FA_cout_986,FA_out_986}=inp_45[48]+inp_46[47]+inp_47[46];
  assign {FA_cout_987,FA_out_987}=inp_45[51]+inp_46[50]+inp_47[49];
  assign {FA_cout_988,FA_out_988}=inp_45[54]+inp_46[53]+inp_47[52];
  assign {FA_cout_989,FA_out_989}=inp_45[57]+inp_46[56]+inp_47[55];
  assign {FA_cout_990,FA_out_990}=inp_45[60]+inp_46[59]+inp_47[58];
  assign {FA_cout_991,FA_out_991}=inp_45[63]+inp_46[62]+inp_47[61];
  assign {FA_cout_992,FA_out_992}=inp_46[18]+inp_47[17]+inp_48[16];
  assign {FA_cout_993,FA_out_993}=inp_46[21]+inp_47[20]+inp_48[19];
  assign {FA_cout_994,FA_out_994}=inp_46[24]+inp_47[23]+inp_48[22];
  assign {FA_cout_995,FA_out_995}=inp_46[27]+inp_47[26]+inp_48[25];
  assign {FA_cout_996,FA_out_996}=inp_46[30]+inp_47[29]+inp_48[28];
  assign {FA_cout_997,FA_out_997}=inp_46[33]+inp_47[32]+inp_48[31];
  assign {FA_cout_998,FA_out_998}=inp_46[36]+inp_47[35]+inp_48[34];
  assign {FA_cout_999,FA_out_999}=inp_46[39]+inp_47[38]+inp_48[37];
  assign {FA_cout_1000,FA_out_1000}=inp_46[42]+inp_47[41]+inp_48[40];
  assign {FA_cout_1001,FA_out_1001}=inp_46[45]+inp_47[44]+inp_48[43];
  assign {FA_cout_1002,FA_out_1002}=inp_46[48]+inp_47[47]+inp_48[46];
  assign {FA_cout_1003,FA_out_1003}=inp_46[51]+inp_47[50]+inp_48[49];
  assign {FA_cout_1004,FA_out_1004}=inp_46[54]+inp_47[53]+inp_48[52];
  assign {FA_cout_1005,FA_out_1005}=inp_46[57]+inp_47[56]+inp_48[55];
  assign {FA_cout_1006,FA_out_1006}=inp_46[60]+inp_47[59]+inp_48[58];
  assign {FA_cout_1007,FA_out_1007}=inp_46[63]+inp_47[62]+inp_48[61];
  assign {FA_cout_1008,FA_out_1008}=inp_47[18]+inp_48[17]+inp_49[16];
  assign {FA_cout_1009,FA_out_1009}=inp_47[21]+inp_48[20]+inp_49[19];
  assign {FA_cout_1010,FA_out_1010}=inp_47[24]+inp_48[23]+inp_49[22];
  assign {FA_cout_1011,FA_out_1011}=inp_47[27]+inp_48[26]+inp_49[25];
  assign {FA_cout_1012,FA_out_1012}=inp_47[30]+inp_48[29]+inp_49[28];
  assign {FA_cout_1013,FA_out_1013}=inp_47[33]+inp_48[32]+inp_49[31];
  assign {FA_cout_1014,FA_out_1014}=inp_47[36]+inp_48[35]+inp_49[34];
  assign {FA_cout_1015,FA_out_1015}=inp_47[39]+inp_48[38]+inp_49[37];
  assign {FA_cout_1016,FA_out_1016}=inp_47[42]+inp_48[41]+inp_49[40];
  assign {FA_cout_1017,FA_out_1017}=inp_47[45]+inp_48[44]+inp_49[43];
  assign {FA_cout_1018,FA_out_1018}=inp_47[48]+inp_48[47]+inp_49[46];
  assign {FA_cout_1019,FA_out_1019}=inp_47[51]+inp_48[50]+inp_49[49];
  assign {FA_cout_1020,FA_out_1020}=inp_47[54]+inp_48[53]+inp_49[52];
  assign {FA_cout_1021,FA_out_1021}=inp_47[57]+inp_48[56]+inp_49[55];
  assign {FA_cout_1022,FA_out_1022}=inp_47[60]+inp_48[59]+inp_49[58];
  assign {FA_cout_1023,FA_out_1023}=inp_47[63]+inp_48[62]+inp_49[61];
  assign {FA_cout_1024,FA_out_1024}=inp_48[2]+inp_49[1]+inp_50[0];
  assign {FA_cout_1025,FA_out_1025}=inp_48[3]+inp_49[2]+inp_50[1];
  assign {FA_cout_1026,FA_out_1026}=inp_48[4]+inp_49[3]+inp_50[2];
  assign {FA_cout_1027,FA_out_1027}=inp_48[5]+inp_49[4]+inp_50[3];
  assign {FA_cout_1028,FA_out_1028}=inp_48[6]+inp_49[5]+inp_50[4];
  assign {FA_cout_1029,FA_out_1029}=inp_48[7]+inp_49[6]+inp_50[5];
  assign {FA_cout_1030,FA_out_1030}=inp_48[8]+inp_49[7]+inp_50[6];
  assign {FA_cout_1031,FA_out_1031}=inp_48[9]+inp_49[8]+inp_50[7];
  assign {FA_cout_1032,FA_out_1032}=inp_48[10]+inp_49[9]+inp_50[8];
  assign {FA_cout_1033,FA_out_1033}=inp_48[11]+inp_49[10]+inp_50[9];
  assign {FA_cout_1034,FA_out_1034}=inp_48[12]+inp_49[11]+inp_50[10];
  assign {FA_cout_1035,FA_out_1035}=inp_48[13]+inp_49[12]+inp_50[11];
  assign {FA_cout_1036,FA_out_1036}=inp_48[14]+inp_49[13]+inp_50[12];
  assign {FA_cout_1037,FA_out_1037}=inp_48[15]+inp_49[14]+inp_50[13];
  assign {FA_cout_1038,FA_out_1038}=inp_48[18]+inp_49[17]+inp_50[16];
  assign {FA_cout_1039,FA_out_1039}=inp_48[21]+inp_49[20]+inp_50[19];
  assign {FA_cout_1040,FA_out_1040}=inp_48[24]+inp_49[23]+inp_50[22];
  assign {FA_cout_1041,FA_out_1041}=inp_48[27]+inp_49[26]+inp_50[25];
  assign {FA_cout_1042,FA_out_1042}=inp_48[30]+inp_49[29]+inp_50[28];
  assign {FA_cout_1043,FA_out_1043}=inp_48[33]+inp_49[32]+inp_50[31];
  assign {FA_cout_1044,FA_out_1044}=inp_48[36]+inp_49[35]+inp_50[34];
  assign {FA_cout_1045,FA_out_1045}=inp_48[39]+inp_49[38]+inp_50[37];
  assign {FA_cout_1046,FA_out_1046}=inp_48[42]+inp_49[41]+inp_50[40];
  assign {FA_cout_1047,FA_out_1047}=inp_48[45]+inp_49[44]+inp_50[43];
  assign {FA_cout_1048,FA_out_1048}=inp_48[48]+inp_49[47]+inp_50[46];
  assign {FA_cout_1049,FA_out_1049}=inp_48[51]+inp_49[50]+inp_50[49];
  assign {FA_cout_1050,FA_out_1050}=inp_48[54]+inp_49[53]+inp_50[52];
  assign {FA_cout_1051,FA_out_1051}=inp_48[57]+inp_49[56]+inp_50[55];
  assign {FA_cout_1052,FA_out_1052}=inp_48[60]+inp_49[59]+inp_50[58];
  assign {FA_cout_1053,FA_out_1053}=inp_48[63]+inp_49[62]+inp_50[61];
  assign {FA_cout_1054,FA_out_1054}=inp_49[15]+inp_50[14]+inp_51[13];
  assign {FA_cout_1055,FA_out_1055}=inp_49[18]+inp_50[17]+inp_51[16];
  assign {FA_cout_1056,FA_out_1056}=inp_49[21]+inp_50[20]+inp_51[19];
  assign {FA_cout_1057,FA_out_1057}=inp_49[24]+inp_50[23]+inp_51[22];
  assign {FA_cout_1058,FA_out_1058}=inp_49[27]+inp_50[26]+inp_51[25];
  assign {FA_cout_1059,FA_out_1059}=inp_49[30]+inp_50[29]+inp_51[28];
  assign {FA_cout_1060,FA_out_1060}=inp_49[33]+inp_50[32]+inp_51[31];
  assign {FA_cout_1061,FA_out_1061}=inp_49[36]+inp_50[35]+inp_51[34];
  assign {FA_cout_1062,FA_out_1062}=inp_49[39]+inp_50[38]+inp_51[37];
  assign {FA_cout_1063,FA_out_1063}=inp_49[42]+inp_50[41]+inp_51[40];
  assign {FA_cout_1064,FA_out_1064}=inp_49[45]+inp_50[44]+inp_51[43];
  assign {FA_cout_1065,FA_out_1065}=inp_49[48]+inp_50[47]+inp_51[46];
  assign {FA_cout_1066,FA_out_1066}=inp_49[51]+inp_50[50]+inp_51[49];
  assign {FA_cout_1067,FA_out_1067}=inp_49[54]+inp_50[53]+inp_51[52];
  assign {FA_cout_1068,FA_out_1068}=inp_49[57]+inp_50[56]+inp_51[55];
  assign {FA_cout_1069,FA_out_1069}=inp_49[60]+inp_50[59]+inp_51[58];
  assign {FA_cout_1070,FA_out_1070}=inp_49[63]+inp_50[62]+inp_51[61];
  assign {FA_cout_1071,FA_out_1071}=inp_50[15]+inp_51[14]+inp_52[13];
  assign {FA_cout_1072,FA_out_1072}=inp_50[18]+inp_51[17]+inp_52[16];
  assign {FA_cout_1073,FA_out_1073}=inp_50[21]+inp_51[20]+inp_52[19];
  assign {FA_cout_1074,FA_out_1074}=inp_50[24]+inp_51[23]+inp_52[22];
  assign {FA_cout_1075,FA_out_1075}=inp_50[27]+inp_51[26]+inp_52[25];
  assign {FA_cout_1076,FA_out_1076}=inp_50[30]+inp_51[29]+inp_52[28];
  assign {FA_cout_1077,FA_out_1077}=inp_50[33]+inp_51[32]+inp_52[31];
  assign {FA_cout_1078,FA_out_1078}=inp_50[36]+inp_51[35]+inp_52[34];
  assign {FA_cout_1079,FA_out_1079}=inp_50[39]+inp_51[38]+inp_52[37];
  assign {FA_cout_1080,FA_out_1080}=inp_50[42]+inp_51[41]+inp_52[40];
  assign {FA_cout_1081,FA_out_1081}=inp_50[45]+inp_51[44]+inp_52[43];
  assign {FA_cout_1082,FA_out_1082}=inp_50[48]+inp_51[47]+inp_52[46];
  assign {FA_cout_1083,FA_out_1083}=inp_50[51]+inp_51[50]+inp_52[49];
  assign {FA_cout_1084,FA_out_1084}=inp_50[54]+inp_51[53]+inp_52[52];
  assign {FA_cout_1085,FA_out_1085}=inp_50[57]+inp_51[56]+inp_52[55];
  assign {FA_cout_1086,FA_out_1086}=inp_50[60]+inp_51[59]+inp_52[58];
  assign {FA_cout_1087,FA_out_1087}=inp_50[63]+inp_51[62]+inp_52[61];
  assign {FA_cout_1088,FA_out_1088}=inp_51[2]+inp_52[1]+inp_53[0];
  assign {FA_cout_1089,FA_out_1089}=inp_51[3]+inp_52[2]+inp_53[1];
  assign {FA_cout_1090,FA_out_1090}=inp_51[4]+inp_52[3]+inp_53[2];
  assign {FA_cout_1091,FA_out_1091}=inp_51[5]+inp_52[4]+inp_53[3];
  assign {FA_cout_1092,FA_out_1092}=inp_51[6]+inp_52[5]+inp_53[4];
  assign {FA_cout_1093,FA_out_1093}=inp_51[7]+inp_52[6]+inp_53[5];
  assign {FA_cout_1094,FA_out_1094}=inp_51[8]+inp_52[7]+inp_53[6];
  assign {FA_cout_1095,FA_out_1095}=inp_51[9]+inp_52[8]+inp_53[7];
  assign {FA_cout_1096,FA_out_1096}=inp_51[10]+inp_52[9]+inp_53[8];
  assign {FA_cout_1097,FA_out_1097}=inp_51[11]+inp_52[10]+inp_53[9];
  assign {FA_cout_1098,FA_out_1098}=inp_51[12]+inp_52[11]+inp_53[10];
  assign {FA_cout_1099,FA_out_1099}=inp_51[15]+inp_52[14]+inp_53[13];
  assign {FA_cout_1100,FA_out_1100}=inp_51[18]+inp_52[17]+inp_53[16];
  assign {FA_cout_1101,FA_out_1101}=inp_51[21]+inp_52[20]+inp_53[19];
  assign {FA_cout_1102,FA_out_1102}=inp_51[24]+inp_52[23]+inp_53[22];
  assign {FA_cout_1103,FA_out_1103}=inp_51[27]+inp_52[26]+inp_53[25];
  assign {FA_cout_1104,FA_out_1104}=inp_51[30]+inp_52[29]+inp_53[28];
  assign {FA_cout_1105,FA_out_1105}=inp_51[33]+inp_52[32]+inp_53[31];
  assign {FA_cout_1106,FA_out_1106}=inp_51[36]+inp_52[35]+inp_53[34];
  assign {FA_cout_1107,FA_out_1107}=inp_51[39]+inp_52[38]+inp_53[37];
  assign {FA_cout_1108,FA_out_1108}=inp_51[42]+inp_52[41]+inp_53[40];
  assign {FA_cout_1109,FA_out_1109}=inp_51[45]+inp_52[44]+inp_53[43];
  assign {FA_cout_1110,FA_out_1110}=inp_51[48]+inp_52[47]+inp_53[46];
  assign {FA_cout_1111,FA_out_1111}=inp_51[51]+inp_52[50]+inp_53[49];
  assign {FA_cout_1112,FA_out_1112}=inp_51[54]+inp_52[53]+inp_53[52];
  assign {FA_cout_1113,FA_out_1113}=inp_51[57]+inp_52[56]+inp_53[55];
  assign {FA_cout_1114,FA_out_1114}=inp_51[60]+inp_52[59]+inp_53[58];
  assign {FA_cout_1115,FA_out_1115}=inp_51[63]+inp_52[62]+inp_53[61];
  assign {FA_cout_1116,FA_out_1116}=inp_52[12]+inp_53[11]+inp_54[10];
  assign {FA_cout_1117,FA_out_1117}=inp_52[15]+inp_53[14]+inp_54[13];
  assign {FA_cout_1118,FA_out_1118}=inp_52[18]+inp_53[17]+inp_54[16];
  assign {FA_cout_1119,FA_out_1119}=inp_52[21]+inp_53[20]+inp_54[19];
  assign {FA_cout_1120,FA_out_1120}=inp_52[24]+inp_53[23]+inp_54[22];
  assign {FA_cout_1121,FA_out_1121}=inp_52[27]+inp_53[26]+inp_54[25];
  assign {FA_cout_1122,FA_out_1122}=inp_52[30]+inp_53[29]+inp_54[28];
  assign {FA_cout_1123,FA_out_1123}=inp_52[33]+inp_53[32]+inp_54[31];
  assign {FA_cout_1124,FA_out_1124}=inp_52[36]+inp_53[35]+inp_54[34];
  assign {FA_cout_1125,FA_out_1125}=inp_52[39]+inp_53[38]+inp_54[37];
  assign {FA_cout_1126,FA_out_1126}=inp_52[42]+inp_53[41]+inp_54[40];
  assign {FA_cout_1127,FA_out_1127}=inp_52[45]+inp_53[44]+inp_54[43];
  assign {FA_cout_1128,FA_out_1128}=inp_52[48]+inp_53[47]+inp_54[46];
  assign {FA_cout_1129,FA_out_1129}=inp_52[51]+inp_53[50]+inp_54[49];
  assign {FA_cout_1130,FA_out_1130}=inp_52[54]+inp_53[53]+inp_54[52];
  assign {FA_cout_1131,FA_out_1131}=inp_52[57]+inp_53[56]+inp_54[55];
  assign {FA_cout_1132,FA_out_1132}=inp_52[60]+inp_53[59]+inp_54[58];
  assign {FA_cout_1133,FA_out_1133}=inp_52[63]+inp_53[62]+inp_54[61];
  assign {FA_cout_1134,FA_out_1134}=inp_53[12]+inp_54[11]+inp_55[10];
  assign {FA_cout_1135,FA_out_1135}=inp_53[15]+inp_54[14]+inp_55[13];
  assign {FA_cout_1136,FA_out_1136}=inp_53[18]+inp_54[17]+inp_55[16];
  assign {FA_cout_1137,FA_out_1137}=inp_53[21]+inp_54[20]+inp_55[19];
  assign {FA_cout_1138,FA_out_1138}=inp_53[24]+inp_54[23]+inp_55[22];
  assign {FA_cout_1139,FA_out_1139}=inp_53[27]+inp_54[26]+inp_55[25];
  assign {FA_cout_1140,FA_out_1140}=inp_53[30]+inp_54[29]+inp_55[28];
  assign {FA_cout_1141,FA_out_1141}=inp_53[33]+inp_54[32]+inp_55[31];
  assign {FA_cout_1142,FA_out_1142}=inp_53[36]+inp_54[35]+inp_55[34];
  assign {FA_cout_1143,FA_out_1143}=inp_53[39]+inp_54[38]+inp_55[37];
  assign {FA_cout_1144,FA_out_1144}=inp_53[42]+inp_54[41]+inp_55[40];
  assign {FA_cout_1145,FA_out_1145}=inp_53[45]+inp_54[44]+inp_55[43];
  assign {FA_cout_1146,FA_out_1146}=inp_53[48]+inp_54[47]+inp_55[46];
  assign {FA_cout_1147,FA_out_1147}=inp_53[51]+inp_54[50]+inp_55[49];
  assign {FA_cout_1148,FA_out_1148}=inp_53[54]+inp_54[53]+inp_55[52];
  assign {FA_cout_1149,FA_out_1149}=inp_53[57]+inp_54[56]+inp_55[55];
  assign {FA_cout_1150,FA_out_1150}=inp_53[60]+inp_54[59]+inp_55[58];
  assign {FA_cout_1151,FA_out_1151}=inp_53[63]+inp_54[62]+inp_55[61];
  assign {FA_cout_1152,FA_out_1152}=inp_54[2]+inp_55[1]+inp_56[0];
  assign {FA_cout_1153,FA_out_1153}=inp_54[3]+inp_55[2]+inp_56[1];
  assign {FA_cout_1154,FA_out_1154}=inp_54[4]+inp_55[3]+inp_56[2];
  assign {FA_cout_1155,FA_out_1155}=inp_54[5]+inp_55[4]+inp_56[3];
  assign {FA_cout_1156,FA_out_1156}=inp_54[6]+inp_55[5]+inp_56[4];
  assign {FA_cout_1157,FA_out_1157}=inp_54[7]+inp_55[6]+inp_56[5];
  assign {FA_cout_1158,FA_out_1158}=inp_54[8]+inp_55[7]+inp_56[6];
  assign {FA_cout_1159,FA_out_1159}=inp_54[9]+inp_55[8]+inp_56[7];
  assign {FA_cout_1160,FA_out_1160}=inp_54[12]+inp_55[11]+inp_56[10];
  assign {FA_cout_1161,FA_out_1161}=inp_54[15]+inp_55[14]+inp_56[13];
  assign {FA_cout_1162,FA_out_1162}=inp_54[18]+inp_55[17]+inp_56[16];
  assign {FA_cout_1163,FA_out_1163}=inp_54[21]+inp_55[20]+inp_56[19];
  assign {FA_cout_1164,FA_out_1164}=inp_54[24]+inp_55[23]+inp_56[22];
  assign {FA_cout_1165,FA_out_1165}=inp_54[27]+inp_55[26]+inp_56[25];
  assign {FA_cout_1166,FA_out_1166}=inp_54[30]+inp_55[29]+inp_56[28];
  assign {FA_cout_1167,FA_out_1167}=inp_54[33]+inp_55[32]+inp_56[31];
  assign {FA_cout_1168,FA_out_1168}=inp_54[36]+inp_55[35]+inp_56[34];
  assign {FA_cout_1169,FA_out_1169}=inp_54[39]+inp_55[38]+inp_56[37];
  assign {FA_cout_1170,FA_out_1170}=inp_54[42]+inp_55[41]+inp_56[40];
  assign {FA_cout_1171,FA_out_1171}=inp_54[45]+inp_55[44]+inp_56[43];
  assign {FA_cout_1172,FA_out_1172}=inp_54[48]+inp_55[47]+inp_56[46];
  assign {FA_cout_1173,FA_out_1173}=inp_54[51]+inp_55[50]+inp_56[49];
  assign {FA_cout_1174,FA_out_1174}=inp_54[54]+inp_55[53]+inp_56[52];
  assign {FA_cout_1175,FA_out_1175}=inp_54[57]+inp_55[56]+inp_56[55];
  assign {FA_cout_1176,FA_out_1176}=inp_54[60]+inp_55[59]+inp_56[58];
  assign {FA_cout_1177,FA_out_1177}=inp_54[63]+inp_55[62]+inp_56[61];
  assign {FA_cout_1178,FA_out_1178}=inp_55[9]+inp_56[8]+inp_57[7];
  assign {FA_cout_1179,FA_out_1179}=inp_55[12]+inp_56[11]+inp_57[10];
  assign {FA_cout_1180,FA_out_1180}=inp_55[15]+inp_56[14]+inp_57[13];
  assign {FA_cout_1181,FA_out_1181}=inp_55[18]+inp_56[17]+inp_57[16];
  assign {FA_cout_1182,FA_out_1182}=inp_55[21]+inp_56[20]+inp_57[19];
  assign {FA_cout_1183,FA_out_1183}=inp_55[24]+inp_56[23]+inp_57[22];
  assign {FA_cout_1184,FA_out_1184}=inp_55[27]+inp_56[26]+inp_57[25];
  assign {FA_cout_1185,FA_out_1185}=inp_55[30]+inp_56[29]+inp_57[28];
  assign {FA_cout_1186,FA_out_1186}=inp_55[33]+inp_56[32]+inp_57[31];
  assign {FA_cout_1187,FA_out_1187}=inp_55[36]+inp_56[35]+inp_57[34];
  assign {FA_cout_1188,FA_out_1188}=inp_55[39]+inp_56[38]+inp_57[37];
  assign {FA_cout_1189,FA_out_1189}=inp_55[42]+inp_56[41]+inp_57[40];
  assign {FA_cout_1190,FA_out_1190}=inp_55[45]+inp_56[44]+inp_57[43];
  assign {FA_cout_1191,FA_out_1191}=inp_55[48]+inp_56[47]+inp_57[46];
  assign {FA_cout_1192,FA_out_1192}=inp_55[51]+inp_56[50]+inp_57[49];
  assign {FA_cout_1193,FA_out_1193}=inp_55[54]+inp_56[53]+inp_57[52];
  assign {FA_cout_1194,FA_out_1194}=inp_55[57]+inp_56[56]+inp_57[55];
  assign {FA_cout_1195,FA_out_1195}=inp_55[60]+inp_56[59]+inp_57[58];
  assign {FA_cout_1196,FA_out_1196}=inp_55[63]+inp_56[62]+inp_57[61];
  assign {FA_cout_1197,FA_out_1197}=inp_56[9]+inp_57[8]+inp_58[7];
  assign {FA_cout_1198,FA_out_1198}=inp_56[12]+inp_57[11]+inp_58[10];
  assign {FA_cout_1199,FA_out_1199}=inp_56[15]+inp_57[14]+inp_58[13];
  assign {FA_cout_1200,FA_out_1200}=inp_56[18]+inp_57[17]+inp_58[16];
  assign {FA_cout_1201,FA_out_1201}=inp_56[21]+inp_57[20]+inp_58[19];
  assign {FA_cout_1202,FA_out_1202}=inp_56[24]+inp_57[23]+inp_58[22];
  assign {FA_cout_1203,FA_out_1203}=inp_56[27]+inp_57[26]+inp_58[25];
  assign {FA_cout_1204,FA_out_1204}=inp_56[30]+inp_57[29]+inp_58[28];
  assign {FA_cout_1205,FA_out_1205}=inp_56[33]+inp_57[32]+inp_58[31];
  assign {FA_cout_1206,FA_out_1206}=inp_56[36]+inp_57[35]+inp_58[34];
  assign {FA_cout_1207,FA_out_1207}=inp_56[39]+inp_57[38]+inp_58[37];
  assign {FA_cout_1208,FA_out_1208}=inp_56[42]+inp_57[41]+inp_58[40];
  assign {FA_cout_1209,FA_out_1209}=inp_56[45]+inp_57[44]+inp_58[43];
  assign {FA_cout_1210,FA_out_1210}=inp_56[48]+inp_57[47]+inp_58[46];
  assign {FA_cout_1211,FA_out_1211}=inp_56[51]+inp_57[50]+inp_58[49];
  assign {FA_cout_1212,FA_out_1212}=inp_56[54]+inp_57[53]+inp_58[52];
  assign {FA_cout_1213,FA_out_1213}=inp_56[57]+inp_57[56]+inp_58[55];
  assign {FA_cout_1214,FA_out_1214}=inp_56[60]+inp_57[59]+inp_58[58];
  assign {FA_cout_1215,FA_out_1215}=inp_56[63]+inp_57[62]+inp_58[61];
  assign {FA_cout_1216,FA_out_1216}=inp_57[2]+inp_58[1]+inp_59[0];
  assign {FA_cout_1217,FA_out_1217}=inp_57[3]+inp_58[2]+inp_59[1];
  assign {FA_cout_1218,FA_out_1218}=inp_57[4]+inp_58[3]+inp_59[2];
  assign {FA_cout_1219,FA_out_1219}=inp_57[5]+inp_58[4]+inp_59[3];
  assign {FA_cout_1220,FA_out_1220}=inp_57[6]+inp_58[5]+inp_59[4];
  assign {FA_cout_1221,FA_out_1221}=inp_57[9]+inp_58[8]+inp_59[7];
  assign {FA_cout_1222,FA_out_1222}=inp_57[12]+inp_58[11]+inp_59[10];
  assign {FA_cout_1223,FA_out_1223}=inp_57[15]+inp_58[14]+inp_59[13];
  assign {FA_cout_1224,FA_out_1224}=inp_57[18]+inp_58[17]+inp_59[16];
  assign {FA_cout_1225,FA_out_1225}=inp_57[21]+inp_58[20]+inp_59[19];
  assign {FA_cout_1226,FA_out_1226}=inp_57[24]+inp_58[23]+inp_59[22];
  assign {FA_cout_1227,FA_out_1227}=inp_57[27]+inp_58[26]+inp_59[25];
  assign {FA_cout_1228,FA_out_1228}=inp_57[30]+inp_58[29]+inp_59[28];
  assign {FA_cout_1229,FA_out_1229}=inp_57[33]+inp_58[32]+inp_59[31];
  assign {FA_cout_1230,FA_out_1230}=inp_57[36]+inp_58[35]+inp_59[34];
  assign {FA_cout_1231,FA_out_1231}=inp_57[39]+inp_58[38]+inp_59[37];
  assign {FA_cout_1232,FA_out_1232}=inp_57[42]+inp_58[41]+inp_59[40];
  assign {FA_cout_1233,FA_out_1233}=inp_57[45]+inp_58[44]+inp_59[43];
  assign {FA_cout_1234,FA_out_1234}=inp_57[48]+inp_58[47]+inp_59[46];
  assign {FA_cout_1235,FA_out_1235}=inp_57[51]+inp_58[50]+inp_59[49];
  assign {FA_cout_1236,FA_out_1236}=inp_57[54]+inp_58[53]+inp_59[52];
  assign {FA_cout_1237,FA_out_1237}=inp_57[57]+inp_58[56]+inp_59[55];
  assign {FA_cout_1238,FA_out_1238}=inp_57[60]+inp_58[59]+inp_59[58];
  assign {FA_cout_1239,FA_out_1239}=inp_57[63]+inp_58[62]+inp_59[61];
  assign {FA_cout_1240,FA_out_1240}=inp_58[6]+inp_59[5]+inp_60[4];
  assign {FA_cout_1241,FA_out_1241}=inp_58[9]+inp_59[8]+inp_60[7];
  assign {FA_cout_1242,FA_out_1242}=inp_58[12]+inp_59[11]+inp_60[10];
  assign {FA_cout_1243,FA_out_1243}=inp_58[15]+inp_59[14]+inp_60[13];
  assign {FA_cout_1244,FA_out_1244}=inp_58[18]+inp_59[17]+inp_60[16];
  assign {FA_cout_1245,FA_out_1245}=inp_58[21]+inp_59[20]+inp_60[19];
  assign {FA_cout_1246,FA_out_1246}=inp_58[24]+inp_59[23]+inp_60[22];
  assign {FA_cout_1247,FA_out_1247}=inp_58[27]+inp_59[26]+inp_60[25];
  assign {FA_cout_1248,FA_out_1248}=inp_58[30]+inp_59[29]+inp_60[28];
  assign {FA_cout_1249,FA_out_1249}=inp_58[33]+inp_59[32]+inp_60[31];
  assign {FA_cout_1250,FA_out_1250}=inp_58[36]+inp_59[35]+inp_60[34];
  assign {FA_cout_1251,FA_out_1251}=inp_58[39]+inp_59[38]+inp_60[37];
  assign {FA_cout_1252,FA_out_1252}=inp_58[42]+inp_59[41]+inp_60[40];
  assign {FA_cout_1253,FA_out_1253}=inp_58[45]+inp_59[44]+inp_60[43];
  assign {FA_cout_1254,FA_out_1254}=inp_58[48]+inp_59[47]+inp_60[46];
  assign {FA_cout_1255,FA_out_1255}=inp_58[51]+inp_59[50]+inp_60[49];
  assign {FA_cout_1256,FA_out_1256}=inp_58[54]+inp_59[53]+inp_60[52];
  assign {FA_cout_1257,FA_out_1257}=inp_58[57]+inp_59[56]+inp_60[55];
  assign {FA_cout_1258,FA_out_1258}=inp_58[60]+inp_59[59]+inp_60[58];
  assign {FA_cout_1259,FA_out_1259}=inp_58[63]+inp_59[62]+inp_60[61];
  assign {FA_cout_1260,FA_out_1260}=inp_59[6]+inp_60[5]+inp_61[4];
  assign {FA_cout_1261,FA_out_1261}=inp_59[9]+inp_60[8]+inp_61[7];
  assign {FA_cout_1262,FA_out_1262}=inp_59[12]+inp_60[11]+inp_61[10];
  assign {FA_cout_1263,FA_out_1263}=inp_59[15]+inp_60[14]+inp_61[13];
  assign {FA_cout_1264,FA_out_1264}=inp_59[18]+inp_60[17]+inp_61[16];
  assign {FA_cout_1265,FA_out_1265}=inp_59[21]+inp_60[20]+inp_61[19];
  assign {FA_cout_1266,FA_out_1266}=inp_59[24]+inp_60[23]+inp_61[22];
  assign {FA_cout_1267,FA_out_1267}=inp_59[27]+inp_60[26]+inp_61[25];
  assign {FA_cout_1268,FA_out_1268}=inp_59[30]+inp_60[29]+inp_61[28];
  assign {FA_cout_1269,FA_out_1269}=inp_59[33]+inp_60[32]+inp_61[31];
  assign {FA_cout_1270,FA_out_1270}=inp_59[36]+inp_60[35]+inp_61[34];
  assign {FA_cout_1271,FA_out_1271}=inp_59[39]+inp_60[38]+inp_61[37];
  assign {FA_cout_1272,FA_out_1272}=inp_59[42]+inp_60[41]+inp_61[40];
  assign {FA_cout_1273,FA_out_1273}=inp_59[45]+inp_60[44]+inp_61[43];
  assign {FA_cout_1274,FA_out_1274}=inp_59[48]+inp_60[47]+inp_61[46];
  assign {FA_cout_1275,FA_out_1275}=inp_59[51]+inp_60[50]+inp_61[49];
  assign {FA_cout_1276,FA_out_1276}=inp_59[54]+inp_60[53]+inp_61[52];
  assign {FA_cout_1277,FA_out_1277}=inp_59[57]+inp_60[56]+inp_61[55];
  assign {FA_cout_1278,FA_out_1278}=inp_59[60]+inp_60[59]+inp_61[58];
  assign {FA_cout_1279,FA_out_1279}=inp_59[63]+inp_60[62]+inp_61[61];
  assign {FA_cout_1280,FA_out_1280}=inp_60[2]+inp_61[1]+inp_62[0];
  assign {FA_cout_1281,FA_out_1281}=inp_60[3]+inp_61[2]+inp_62[1];
  assign {FA_cout_1282,FA_out_1282}=inp_60[6]+inp_61[5]+inp_62[4];
  assign {FA_cout_1283,FA_out_1283}=inp_60[9]+inp_61[8]+inp_62[7];
  assign {FA_cout_1284,FA_out_1284}=inp_60[12]+inp_61[11]+inp_62[10];
  assign {FA_cout_1285,FA_out_1285}=inp_60[15]+inp_61[14]+inp_62[13];
  assign {FA_cout_1286,FA_out_1286}=inp_60[18]+inp_61[17]+inp_62[16];
  assign {FA_cout_1287,FA_out_1287}=inp_60[21]+inp_61[20]+inp_62[19];
  assign {FA_cout_1288,FA_out_1288}=inp_60[24]+inp_61[23]+inp_62[22];
  assign {FA_cout_1289,FA_out_1289}=inp_60[27]+inp_61[26]+inp_62[25];
  assign {FA_cout_1290,FA_out_1290}=inp_60[30]+inp_61[29]+inp_62[28];
  assign {FA_cout_1291,FA_out_1291}=inp_60[33]+inp_61[32]+inp_62[31];
  assign {FA_cout_1292,FA_out_1292}=inp_60[36]+inp_61[35]+inp_62[34];
  assign {FA_cout_1293,FA_out_1293}=inp_60[39]+inp_61[38]+inp_62[37];
  assign {FA_cout_1294,FA_out_1294}=inp_60[42]+inp_61[41]+inp_62[40];
  assign {FA_cout_1295,FA_out_1295}=inp_60[45]+inp_61[44]+inp_62[43];
  assign {FA_cout_1296,FA_out_1296}=inp_60[48]+inp_61[47]+inp_62[46];
  assign {FA_cout_1297,FA_out_1297}=inp_60[51]+inp_61[50]+inp_62[49];
  assign {FA_cout_1298,FA_out_1298}=inp_60[54]+inp_61[53]+inp_62[52];
  assign {FA_cout_1299,FA_out_1299}=inp_60[57]+inp_61[56]+inp_62[55];
  assign {FA_cout_1300,FA_out_1300}=inp_60[60]+inp_61[59]+inp_62[58];
  assign {FA_cout_1301,FA_out_1301}=inp_60[63]+inp_61[62]+inp_62[61];
  assign {FA_cout_1302,FA_out_1302}=inp_61[3]+inp_62[2]+inp_63[1];
  assign {FA_cout_1303,FA_out_1303}=inp_61[6]+inp_62[5]+inp_63[4];
  assign {FA_cout_1304,FA_out_1304}=inp_61[9]+inp_62[8]+inp_63[7];
  assign {FA_cout_1305,FA_out_1305}=inp_61[12]+inp_62[11]+inp_63[10];
  assign {FA_cout_1306,FA_out_1306}=inp_61[15]+inp_62[14]+inp_63[13];
  assign {FA_cout_1307,FA_out_1307}=inp_61[18]+inp_62[17]+inp_63[16];
  assign {FA_cout_1308,FA_out_1308}=inp_61[21]+inp_62[20]+inp_63[19];
  assign {FA_cout_1309,FA_out_1309}=inp_61[24]+inp_62[23]+inp_63[22];
  assign {FA_cout_1310,FA_out_1310}=inp_61[27]+inp_62[26]+inp_63[25];
  assign {FA_cout_1311,FA_out_1311}=inp_61[30]+inp_62[29]+inp_63[28];
  assign {FA_cout_1312,FA_out_1312}=inp_61[33]+inp_62[32]+inp_63[31];
  assign {FA_cout_1313,FA_out_1313}=inp_61[36]+inp_62[35]+inp_63[34];
  assign {FA_cout_1314,FA_out_1314}=inp_61[39]+inp_62[38]+inp_63[37];
  assign {FA_cout_1315,FA_out_1315}=inp_61[42]+inp_62[41]+inp_63[40];
  assign {FA_cout_1316,FA_out_1316}=inp_61[45]+inp_62[44]+inp_63[43];
  assign {FA_cout_1317,FA_out_1317}=inp_61[48]+inp_62[47]+inp_63[46];
  assign {FA_cout_1318,FA_out_1318}=inp_61[51]+inp_62[50]+inp_63[49];
  assign {FA_cout_1319,FA_out_1319}=inp_61[54]+inp_62[53]+inp_63[52];
  assign {FA_cout_1320,FA_out_1320}=inp_61[57]+inp_62[56]+inp_63[55];
  assign {FA_cout_1321,FA_out_1321}=inp_61[60]+inp_62[59]+inp_63[58];
  assign {FA_cout_1322,FA_out_1322}=inp_61[63]+inp_62[62]+inp_63[61];
  assign {FA_cout_1323,FA_out_1323}=FA_cout_0+FA_out_1+inp_3[0];
  assign {FA_cout_1324,FA_out_1324}=FA_cout_1+FA_out_2+HA_out_1;
  assign {FA_cout_1325,FA_out_1325}=FA_cout_2+FA_out_3+HA_cout_1;
  assign {FA_cout_1326,FA_out_1326}=FA_cout_3+FA_out_4+FA_cout_64;
  assign {FA_cout_1327,FA_out_1327}=FA_cout_4+FA_out_5+FA_cout_65;
  assign {FA_cout_1328,FA_out_1328}=FA_cout_5+FA_out_6+FA_cout_66;
  assign {FA_cout_1329,FA_out_1329}=FA_cout_6+FA_out_7+FA_cout_67;
  assign {FA_cout_1330,FA_out_1330}=FA_cout_7+FA_out_8+FA_cout_68;
  assign {FA_cout_1331,FA_out_1331}=FA_cout_8+FA_out_9+FA_cout_69;
  assign {FA_cout_1332,FA_out_1332}=FA_cout_9+FA_out_10+FA_cout_70;
  assign {FA_cout_1333,FA_out_1333}=FA_cout_10+FA_out_11+FA_cout_71;
  assign {FA_cout_1334,FA_out_1334}=FA_cout_11+FA_out_12+FA_cout_72;
  assign {FA_cout_1335,FA_out_1335}=FA_cout_12+FA_out_13+FA_cout_73;
  assign {FA_cout_1336,FA_out_1336}=FA_cout_13+FA_out_14+FA_cout_74;
  assign {FA_cout_1337,FA_out_1337}=FA_cout_14+FA_out_15+FA_cout_75;
  assign {FA_cout_1338,FA_out_1338}=FA_cout_15+FA_out_16+FA_cout_76;
  assign {FA_cout_1339,FA_out_1339}=FA_cout_16+FA_out_17+FA_cout_77;
  assign {FA_cout_1340,FA_out_1340}=FA_cout_17+FA_out_18+FA_cout_78;
  assign {FA_cout_1341,FA_out_1341}=FA_cout_18+FA_out_19+FA_cout_79;
  assign {FA_cout_1342,FA_out_1342}=FA_cout_19+FA_out_20+FA_cout_80;
  assign {FA_cout_1343,FA_out_1343}=FA_cout_20+FA_out_21+FA_cout_81;
  assign {FA_cout_1344,FA_out_1344}=FA_cout_21+FA_out_22+FA_cout_82;
  assign {FA_cout_1345,FA_out_1345}=FA_cout_22+FA_out_23+FA_cout_83;
  assign {FA_cout_1346,FA_out_1346}=FA_cout_23+FA_out_24+FA_cout_84;
  assign {FA_cout_1347,FA_out_1347}=FA_cout_24+FA_out_25+FA_cout_85;
  assign {FA_cout_1348,FA_out_1348}=FA_cout_25+FA_out_26+FA_cout_86;
  assign {FA_cout_1349,FA_out_1349}=FA_cout_26+FA_out_27+FA_cout_87;
  assign {FA_cout_1350,FA_out_1350}=FA_cout_27+FA_out_28+FA_cout_88;
  assign {FA_cout_1351,FA_out_1351}=FA_cout_28+FA_out_29+FA_cout_89;
  assign {FA_cout_1352,FA_out_1352}=FA_cout_29+FA_out_30+FA_cout_90;
  assign {FA_cout_1353,FA_out_1353}=FA_cout_30+FA_out_31+FA_cout_91;
  assign {FA_cout_1354,FA_out_1354}=FA_cout_31+FA_out_32+FA_cout_92;
  assign {FA_cout_1355,FA_out_1355}=FA_cout_32+FA_out_33+FA_cout_93;
  assign {FA_cout_1356,FA_out_1356}=FA_cout_33+FA_out_34+FA_cout_94;
  assign {FA_cout_1357,FA_out_1357}=FA_cout_34+FA_out_35+FA_cout_95;
  assign {FA_cout_1358,FA_out_1358}=FA_cout_35+FA_out_36+FA_cout_96;
  assign {FA_cout_1359,FA_out_1359}=FA_cout_36+FA_out_37+FA_cout_97;
  assign {FA_cout_1360,FA_out_1360}=FA_cout_37+FA_out_38+FA_cout_98;
  assign {FA_cout_1361,FA_out_1361}=FA_cout_38+FA_out_39+FA_cout_99;
  assign {FA_cout_1362,FA_out_1362}=FA_cout_39+FA_out_40+FA_cout_100;
  assign {FA_cout_1363,FA_out_1363}=FA_cout_40+FA_out_41+FA_cout_101;
  assign {FA_cout_1364,FA_out_1364}=FA_cout_41+FA_out_42+FA_cout_102;
  assign {FA_cout_1365,FA_out_1365}=FA_cout_42+FA_out_43+FA_cout_103;
  assign {FA_cout_1366,FA_out_1366}=FA_cout_43+FA_out_44+FA_cout_104;
  assign {FA_cout_1367,FA_out_1367}=FA_cout_44+FA_out_45+FA_cout_105;
  assign {FA_cout_1368,FA_out_1368}=FA_cout_45+FA_out_46+FA_cout_106;
  assign {FA_cout_1369,FA_out_1369}=FA_cout_46+FA_out_47+FA_cout_107;
  assign {FA_cout_1370,FA_out_1370}=FA_cout_47+FA_out_48+FA_cout_108;
  assign {FA_cout_1371,FA_out_1371}=FA_cout_48+FA_out_49+FA_cout_109;
  assign {FA_cout_1372,FA_out_1372}=FA_cout_49+FA_out_50+FA_cout_110;
  assign {FA_cout_1373,FA_out_1373}=FA_cout_50+FA_out_51+FA_cout_111;
  assign {FA_cout_1374,FA_out_1374}=FA_cout_51+FA_out_52+FA_cout_112;
  assign {FA_cout_1375,FA_out_1375}=FA_cout_52+FA_out_53+FA_cout_113;
  assign {FA_cout_1376,FA_out_1376}=FA_cout_53+FA_out_54+FA_cout_114;
  assign {FA_cout_1377,FA_out_1377}=FA_cout_54+FA_out_55+FA_cout_115;
  assign {FA_cout_1378,FA_out_1378}=FA_cout_55+FA_out_56+FA_cout_116;
  assign {FA_cout_1379,FA_out_1379}=FA_cout_56+FA_out_57+FA_cout_117;
  assign {FA_cout_1380,FA_out_1380}=FA_cout_57+FA_out_58+FA_cout_118;
  assign {FA_cout_1381,FA_out_1381}=FA_cout_58+FA_out_59+FA_cout_119;
  assign {FA_cout_1382,FA_out_1382}=FA_cout_59+FA_out_60+FA_cout_120;
  assign {FA_cout_1383,FA_out_1383}=FA_cout_60+FA_out_61+FA_cout_121;
  assign {FA_cout_1384,FA_out_1384}=FA_cout_61+FA_out_62+FA_cout_122;
  assign {FA_cout_1385,FA_out_1385}=FA_cout_62+FA_out_63+FA_cout_124;
  assign {FA_cout_1386,FA_out_1386}=FA_cout_63+FA_out_123+FA_cout_126;
  assign {FA_cout_1387,FA_out_1387}=FA_cout_123+FA_out_125+FA_cout_184;
  assign {FA_cout_1388,FA_out_1388}=FA_out_67+HA_cout_2+FA_out_128;
  assign {FA_cout_1389,FA_out_1389}=FA_out_68+FA_cout_128+FA_out_129;
  assign {FA_cout_1390,FA_out_1390}=FA_out_69+FA_cout_129+FA_out_130;
  assign {FA_cout_1391,FA_out_1391}=FA_out_70+FA_cout_130+FA_out_131;
  assign {FA_cout_1392,FA_out_1392}=FA_out_71+FA_cout_131+FA_out_132;
  assign {FA_cout_1393,FA_out_1393}=FA_out_72+FA_cout_132+FA_out_133;
  assign {FA_cout_1394,FA_out_1394}=FA_out_73+FA_cout_133+FA_out_134;
  assign {FA_cout_1395,FA_out_1395}=FA_out_74+FA_cout_134+FA_out_135;
  assign {FA_cout_1396,FA_out_1396}=FA_out_75+FA_cout_135+FA_out_136;
  assign {FA_cout_1397,FA_out_1397}=FA_out_76+FA_cout_136+FA_out_137;
  assign {FA_cout_1398,FA_out_1398}=FA_out_77+FA_cout_137+FA_out_138;
  assign {FA_cout_1399,FA_out_1399}=FA_out_78+FA_cout_138+FA_out_139;
  assign {FA_cout_1400,FA_out_1400}=FA_out_79+FA_cout_139+FA_out_140;
  assign {FA_cout_1401,FA_out_1401}=FA_out_80+FA_cout_140+FA_out_141;
  assign {FA_cout_1402,FA_out_1402}=FA_out_81+FA_cout_141+FA_out_142;
  assign {FA_cout_1403,FA_out_1403}=FA_out_82+FA_cout_142+FA_out_143;
  assign {FA_cout_1404,FA_out_1404}=FA_out_83+FA_cout_143+FA_out_144;
  assign {FA_cout_1405,FA_out_1405}=FA_out_84+FA_cout_144+FA_out_145;
  assign {FA_cout_1406,FA_out_1406}=FA_out_85+FA_cout_145+FA_out_146;
  assign {FA_cout_1407,FA_out_1407}=FA_out_86+FA_cout_146+FA_out_147;
  assign {FA_cout_1408,FA_out_1408}=FA_out_87+FA_cout_147+FA_out_148;
  assign {FA_cout_1409,FA_out_1409}=FA_out_88+FA_cout_148+FA_out_149;
  assign {FA_cout_1410,FA_out_1410}=FA_out_89+FA_cout_149+FA_out_150;
  assign {FA_cout_1411,FA_out_1411}=FA_out_90+FA_cout_150+FA_out_151;
  assign {FA_cout_1412,FA_out_1412}=FA_out_91+FA_cout_151+FA_out_152;
  assign {FA_cout_1413,FA_out_1413}=FA_out_92+FA_cout_152+FA_out_153;
  assign {FA_cout_1414,FA_out_1414}=FA_out_93+FA_cout_153+FA_out_154;
  assign {FA_cout_1415,FA_out_1415}=FA_out_94+FA_cout_154+FA_out_155;
  assign {FA_cout_1416,FA_out_1416}=FA_out_95+FA_cout_155+FA_out_156;
  assign {FA_cout_1417,FA_out_1417}=FA_out_96+FA_cout_156+FA_out_157;
  assign {FA_cout_1418,FA_out_1418}=FA_out_97+FA_cout_157+FA_out_158;
  assign {FA_cout_1419,FA_out_1419}=FA_out_98+FA_cout_158+FA_out_159;
  assign {FA_cout_1420,FA_out_1420}=FA_out_99+FA_cout_159+FA_out_160;
  assign {FA_cout_1421,FA_out_1421}=FA_out_100+FA_cout_160+FA_out_161;
  assign {FA_cout_1422,FA_out_1422}=FA_out_101+FA_cout_161+FA_out_162;
  assign {FA_cout_1423,FA_out_1423}=FA_out_102+FA_cout_162+FA_out_163;
  assign {FA_cout_1424,FA_out_1424}=FA_out_103+FA_cout_163+FA_out_164;
  assign {FA_cout_1425,FA_out_1425}=FA_out_104+FA_cout_164+FA_out_165;
  assign {FA_cout_1426,FA_out_1426}=FA_out_105+FA_cout_165+FA_out_166;
  assign {FA_cout_1427,FA_out_1427}=FA_out_106+FA_cout_166+FA_out_167;
  assign {FA_cout_1428,FA_out_1428}=FA_out_107+FA_cout_167+FA_out_168;
  assign {FA_cout_1429,FA_out_1429}=FA_out_108+FA_cout_168+FA_out_169;
  assign {FA_cout_1430,FA_out_1430}=FA_out_109+FA_cout_169+FA_out_170;
  assign {FA_cout_1431,FA_out_1431}=FA_out_110+FA_cout_170+FA_out_171;
  assign {FA_cout_1432,FA_out_1432}=FA_out_111+FA_cout_171+FA_out_172;
  assign {FA_cout_1433,FA_out_1433}=FA_out_112+FA_cout_172+FA_out_173;
  assign {FA_cout_1434,FA_out_1434}=FA_out_113+FA_cout_173+FA_out_174;
  assign {FA_cout_1435,FA_out_1435}=FA_out_114+FA_cout_174+FA_out_175;
  assign {FA_cout_1436,FA_out_1436}=FA_out_115+FA_cout_175+FA_out_176;
  assign {FA_cout_1437,FA_out_1437}=FA_out_116+FA_cout_176+FA_out_177;
  assign {FA_cout_1438,FA_out_1438}=FA_out_117+FA_cout_177+FA_out_178;
  assign {FA_cout_1439,FA_out_1439}=FA_out_118+FA_cout_178+FA_out_179;
  assign {FA_cout_1440,FA_out_1440}=FA_out_119+FA_cout_179+FA_out_180;
  assign {FA_cout_1441,FA_out_1441}=FA_out_120+FA_cout_180+FA_out_181;
  assign {FA_cout_1442,FA_out_1442}=FA_out_121+FA_cout_181+FA_out_182;
  assign {FA_cout_1443,FA_out_1443}=FA_out_122+FA_cout_182+FA_out_183;
  assign {FA_cout_1444,FA_out_1444}=FA_out_124+FA_cout_183+FA_out_186;
  assign {FA_cout_1445,FA_out_1445}=FA_cout_125+FA_out_127+FA_cout_187;
  assign {FA_cout_1446,FA_out_1446}=FA_out_126+FA_cout_186+FA_out_189;
  assign {FA_cout_1447,FA_out_1447}=FA_cout_127+FA_out_185+FA_cout_190;
  assign {FA_cout_1448,FA_out_1448}=FA_out_184+FA_cout_189+FA_out_245;
  assign {FA_cout_1449,FA_out_1449}=FA_cout_185+FA_out_188+FA_cout_246;
  assign {FA_cout_1450,FA_out_1450}=FA_out_187+FA_cout_245+FA_out_249;
  assign {FA_cout_1451,FA_out_1451}=FA_cout_188+FA_out_191+FA_cout_250;
  assign {FA_cout_1452,FA_out_1452}=FA_out_190+FA_cout_249+FA_out_253;
  assign {FA_cout_1453,FA_out_1453}=FA_cout_191+FA_out_247+FA_cout_254;
  assign {FA_cout_1454,FA_out_1454}=FA_cout_192+FA_out_193+inp_12[0];
  assign {FA_cout_1455,FA_out_1455}=FA_cout_193+FA_out_194+HA_out_4;
  assign {FA_cout_1456,FA_out_1456}=FA_cout_194+FA_out_195+HA_cout_4;
  assign {FA_cout_1457,FA_out_1457}=FA_cout_195+FA_out_196+FA_cout_256;
  assign {FA_cout_1458,FA_out_1458}=FA_cout_196+FA_out_197+FA_cout_257;
  assign {FA_cout_1459,FA_out_1459}=FA_cout_197+FA_out_198+FA_cout_258;
  assign {FA_cout_1460,FA_out_1460}=FA_cout_198+FA_out_199+FA_cout_259;
  assign {FA_cout_1461,FA_out_1461}=FA_cout_199+FA_out_200+FA_cout_260;
  assign {FA_cout_1462,FA_out_1462}=FA_cout_200+FA_out_201+FA_cout_261;
  assign {FA_cout_1463,FA_out_1463}=FA_cout_201+FA_out_202+FA_cout_262;
  assign {FA_cout_1464,FA_out_1464}=FA_cout_202+FA_out_203+FA_cout_263;
  assign {FA_cout_1465,FA_out_1465}=FA_cout_203+FA_out_204+FA_cout_264;
  assign {FA_cout_1466,FA_out_1466}=FA_cout_204+FA_out_205+FA_cout_265;
  assign {FA_cout_1467,FA_out_1467}=FA_cout_205+FA_out_206+FA_cout_266;
  assign {FA_cout_1468,FA_out_1468}=FA_cout_206+FA_out_207+FA_cout_267;
  assign {FA_cout_1469,FA_out_1469}=FA_cout_207+FA_out_208+FA_cout_268;
  assign {FA_cout_1470,FA_out_1470}=FA_cout_208+FA_out_209+FA_cout_269;
  assign {FA_cout_1471,FA_out_1471}=FA_cout_209+FA_out_210+FA_cout_270;
  assign {FA_cout_1472,FA_out_1472}=FA_cout_210+FA_out_211+FA_cout_271;
  assign {FA_cout_1473,FA_out_1473}=FA_cout_211+FA_out_212+FA_cout_272;
  assign {FA_cout_1474,FA_out_1474}=FA_cout_212+FA_out_213+FA_cout_273;
  assign {FA_cout_1475,FA_out_1475}=FA_cout_213+FA_out_214+FA_cout_274;
  assign {FA_cout_1476,FA_out_1476}=FA_cout_214+FA_out_215+FA_cout_275;
  assign {FA_cout_1477,FA_out_1477}=FA_cout_215+FA_out_216+FA_cout_276;
  assign {FA_cout_1478,FA_out_1478}=FA_cout_216+FA_out_217+FA_cout_277;
  assign {FA_cout_1479,FA_out_1479}=FA_cout_217+FA_out_218+FA_cout_278;
  assign {FA_cout_1480,FA_out_1480}=FA_cout_218+FA_out_219+FA_cout_279;
  assign {FA_cout_1481,FA_out_1481}=FA_cout_219+FA_out_220+FA_cout_280;
  assign {FA_cout_1482,FA_out_1482}=FA_cout_220+FA_out_221+FA_cout_281;
  assign {FA_cout_1483,FA_out_1483}=FA_cout_221+FA_out_222+FA_cout_282;
  assign {FA_cout_1484,FA_out_1484}=FA_cout_222+FA_out_223+FA_cout_283;
  assign {FA_cout_1485,FA_out_1485}=FA_cout_223+FA_out_224+FA_cout_284;
  assign {FA_cout_1486,FA_out_1486}=FA_cout_224+FA_out_225+FA_cout_285;
  assign {FA_cout_1487,FA_out_1487}=FA_cout_225+FA_out_226+FA_cout_286;
  assign {FA_cout_1488,FA_out_1488}=FA_cout_226+FA_out_227+FA_cout_287;
  assign {FA_cout_1489,FA_out_1489}=FA_cout_227+FA_out_228+FA_cout_288;
  assign {FA_cout_1490,FA_out_1490}=FA_cout_228+FA_out_229+FA_cout_289;
  assign {FA_cout_1491,FA_out_1491}=FA_cout_229+FA_out_230+FA_cout_290;
  assign {FA_cout_1492,FA_out_1492}=FA_cout_230+FA_out_231+FA_cout_291;
  assign {FA_cout_1493,FA_out_1493}=FA_cout_231+FA_out_232+FA_cout_292;
  assign {FA_cout_1494,FA_out_1494}=FA_cout_232+FA_out_233+FA_cout_293;
  assign {FA_cout_1495,FA_out_1495}=FA_cout_233+FA_out_234+FA_cout_294;
  assign {FA_cout_1496,FA_out_1496}=FA_cout_234+FA_out_235+FA_cout_295;
  assign {FA_cout_1497,FA_out_1497}=FA_cout_235+FA_out_236+FA_cout_296;
  assign {FA_cout_1498,FA_out_1498}=FA_cout_236+FA_out_237+FA_cout_297;
  assign {FA_cout_1499,FA_out_1499}=FA_cout_237+FA_out_238+FA_cout_298;
  assign {FA_cout_1500,FA_out_1500}=FA_cout_238+FA_out_239+FA_cout_299;
  assign {FA_cout_1501,FA_out_1501}=FA_cout_239+FA_out_240+FA_cout_300;
  assign {FA_cout_1502,FA_out_1502}=FA_cout_240+FA_out_241+FA_cout_301;
  assign {FA_cout_1503,FA_out_1503}=FA_cout_241+FA_out_242+FA_cout_302;
  assign {FA_cout_1504,FA_out_1504}=FA_cout_242+FA_out_243+FA_cout_303;
  assign {FA_cout_1505,FA_out_1505}=FA_cout_243+FA_out_244+FA_cout_304;
  assign {FA_cout_1506,FA_out_1506}=FA_cout_244+FA_out_248+FA_cout_305;
  assign {FA_cout_1507,FA_out_1507}=FA_out_246+FA_cout_253+FA_out_307;
  assign {FA_cout_1508,FA_out_1508}=FA_cout_247+FA_out_251+FA_cout_308;
  assign {FA_cout_1509,FA_out_1509}=FA_cout_248+FA_out_252+FA_cout_310;
  assign {FA_cout_1510,FA_out_1510}=FA_out_250+FA_cout_307+FA_out_312;
  assign {FA_cout_1511,FA_out_1511}=FA_cout_251+FA_out_255+FA_cout_313;
  assign {FA_cout_1512,FA_out_1512}=FA_cout_252+FA_out_306+FA_cout_315;
  assign {FA_cout_1513,FA_out_1513}=FA_out_254+FA_cout_312+FA_out_317;
  assign {FA_cout_1514,FA_out_1514}=FA_cout_255+FA_out_309+FA_cout_318;
  assign {FA_cout_1515,FA_out_1515}=FA_cout_306+FA_out_311+FA_cout_367;
  assign {FA_cout_1516,FA_out_1516}=FA_out_308+FA_cout_317+FA_out_369;
  assign {FA_cout_1517,FA_out_1517}=FA_cout_309+FA_out_314+FA_cout_370;
  assign {FA_cout_1518,FA_out_1518}=FA_out_259+HA_cout_5+FA_out_320;
  assign {FA_cout_1519,FA_out_1519}=FA_out_260+FA_cout_320+FA_out_321;
  assign {FA_cout_1520,FA_out_1520}=FA_out_261+FA_cout_321+FA_out_322;
  assign {FA_cout_1521,FA_out_1521}=FA_out_262+FA_cout_322+FA_out_323;
  assign {FA_cout_1522,FA_out_1522}=FA_out_263+FA_cout_323+FA_out_324;
  assign {FA_cout_1523,FA_out_1523}=FA_out_264+FA_cout_324+FA_out_325;
  assign {FA_cout_1524,FA_out_1524}=FA_out_265+FA_cout_325+FA_out_326;
  assign {FA_cout_1525,FA_out_1525}=FA_out_266+FA_cout_326+FA_out_327;
  assign {FA_cout_1526,FA_out_1526}=FA_out_267+FA_cout_327+FA_out_328;
  assign {FA_cout_1527,FA_out_1527}=FA_out_268+FA_cout_328+FA_out_329;
  assign {FA_cout_1528,FA_out_1528}=FA_out_269+FA_cout_329+FA_out_330;
  assign {FA_cout_1529,FA_out_1529}=FA_out_270+FA_cout_330+FA_out_331;
  assign {FA_cout_1530,FA_out_1530}=FA_out_271+FA_cout_331+FA_out_332;
  assign {FA_cout_1531,FA_out_1531}=FA_out_272+FA_cout_332+FA_out_333;
  assign {FA_cout_1532,FA_out_1532}=FA_out_273+FA_cout_333+FA_out_334;
  assign {FA_cout_1533,FA_out_1533}=FA_out_274+FA_cout_334+FA_out_335;
  assign {FA_cout_1534,FA_out_1534}=FA_out_275+FA_cout_335+FA_out_336;
  assign {FA_cout_1535,FA_out_1535}=FA_out_276+FA_cout_336+FA_out_337;
  assign {FA_cout_1536,FA_out_1536}=FA_out_277+FA_cout_337+FA_out_338;
  assign {FA_cout_1537,FA_out_1537}=FA_out_278+FA_cout_338+FA_out_339;
  assign {FA_cout_1538,FA_out_1538}=FA_out_279+FA_cout_339+FA_out_340;
  assign {FA_cout_1539,FA_out_1539}=FA_out_280+FA_cout_340+FA_out_341;
  assign {FA_cout_1540,FA_out_1540}=FA_out_281+FA_cout_341+FA_out_342;
  assign {FA_cout_1541,FA_out_1541}=FA_out_282+FA_cout_342+FA_out_343;
  assign {FA_cout_1542,FA_out_1542}=FA_out_283+FA_cout_343+FA_out_344;
  assign {FA_cout_1543,FA_out_1543}=FA_out_284+FA_cout_344+FA_out_345;
  assign {FA_cout_1544,FA_out_1544}=FA_out_285+FA_cout_345+FA_out_346;
  assign {FA_cout_1545,FA_out_1545}=FA_out_286+FA_cout_346+FA_out_347;
  assign {FA_cout_1546,FA_out_1546}=FA_out_287+FA_cout_347+FA_out_348;
  assign {FA_cout_1547,FA_out_1547}=FA_out_288+FA_cout_348+FA_out_349;
  assign {FA_cout_1548,FA_out_1548}=FA_out_289+FA_cout_349+FA_out_350;
  assign {FA_cout_1549,FA_out_1549}=FA_out_290+FA_cout_350+FA_out_351;
  assign {FA_cout_1550,FA_out_1550}=FA_out_291+FA_cout_351+FA_out_352;
  assign {FA_cout_1551,FA_out_1551}=FA_out_292+FA_cout_352+FA_out_353;
  assign {FA_cout_1552,FA_out_1552}=FA_out_293+FA_cout_353+FA_out_354;
  assign {FA_cout_1553,FA_out_1553}=FA_out_294+FA_cout_354+FA_out_355;
  assign {FA_cout_1554,FA_out_1554}=FA_out_295+FA_cout_355+FA_out_356;
  assign {FA_cout_1555,FA_out_1555}=FA_out_296+FA_cout_356+FA_out_357;
  assign {FA_cout_1556,FA_out_1556}=FA_out_297+FA_cout_357+FA_out_358;
  assign {FA_cout_1557,FA_out_1557}=FA_out_298+FA_cout_358+FA_out_359;
  assign {FA_cout_1558,FA_out_1558}=FA_out_299+FA_cout_359+FA_out_360;
  assign {FA_cout_1559,FA_out_1559}=FA_out_300+FA_cout_360+FA_out_361;
  assign {FA_cout_1560,FA_out_1560}=FA_out_301+FA_cout_361+FA_out_362;
  assign {FA_cout_1561,FA_out_1561}=FA_out_302+FA_cout_362+FA_out_363;
  assign {FA_cout_1562,FA_out_1562}=FA_out_303+FA_cout_363+FA_out_364;
  assign {FA_cout_1563,FA_out_1563}=FA_out_304+FA_cout_364+FA_out_365;
  assign {FA_cout_1564,FA_out_1564}=FA_out_305+FA_cout_365+FA_out_366;
  assign {FA_cout_1565,FA_out_1565}=FA_out_310+FA_cout_366+FA_out_372;
  assign {FA_cout_1566,FA_out_1566}=FA_cout_311+FA_out_316+FA_cout_373;
  assign {FA_cout_1567,FA_out_1567}=FA_out_313+FA_cout_369+FA_out_375;
  assign {FA_cout_1568,FA_out_1568}=FA_cout_314+FA_out_319+FA_cout_376;
  assign {FA_cout_1569,FA_out_1569}=FA_out_315+FA_cout_372+FA_out_378;
  assign {FA_cout_1570,FA_out_1570}=FA_cout_316+FA_out_368+FA_cout_379;
  assign {FA_cout_1571,FA_out_1571}=FA_out_318+FA_cout_375+FA_out_381;
  assign {FA_cout_1572,FA_out_1572}=FA_cout_319+FA_out_371+FA_cout_382;
  assign {FA_cout_1573,FA_out_1573}=FA_out_367+FA_cout_378+FA_out_428;
  assign {FA_cout_1574,FA_out_1574}=FA_cout_368+FA_out_374+FA_cout_429;
  assign {FA_cout_1575,FA_out_1575}=FA_out_370+FA_cout_381+FA_out_431;
  assign {FA_cout_1576,FA_out_1576}=FA_cout_371+FA_out_377+FA_cout_432;
  assign {FA_cout_1577,FA_out_1577}=FA_out_373+FA_cout_428+FA_out_435;
  assign {FA_cout_1578,FA_out_1578}=FA_cout_374+FA_out_380+FA_cout_436;
  assign {FA_cout_1579,FA_out_1579}=FA_out_376+FA_cout_431+FA_out_438;
  assign {FA_cout_1580,FA_out_1580}=FA_cout_377+FA_out_383+FA_cout_439;
  assign {FA_cout_1581,FA_out_1581}=FA_out_379+FA_cout_435+FA_out_442;
  assign {FA_cout_1582,FA_out_1582}=FA_cout_380+FA_out_430+FA_cout_443;
  assign {FA_cout_1583,FA_out_1583}=FA_out_382+FA_cout_438+FA_out_445;
  assign {FA_cout_1584,FA_out_1584}=FA_cout_383+FA_out_433+FA_cout_446;
  assign {FA_cout_1585,FA_out_1585}=FA_cout_384+FA_out_385+inp_21[0];
  assign {FA_cout_1586,FA_out_1586}=FA_cout_385+FA_out_386+HA_out_7;
  assign {FA_cout_1587,FA_out_1587}=FA_cout_386+FA_out_387+HA_cout_7;
  assign {FA_cout_1588,FA_out_1588}=FA_cout_387+FA_out_388+FA_cout_448;
  assign {FA_cout_1589,FA_out_1589}=FA_cout_388+FA_out_389+FA_cout_449;
  assign {FA_cout_1590,FA_out_1590}=FA_cout_389+FA_out_390+FA_cout_450;
  assign {FA_cout_1591,FA_out_1591}=FA_cout_390+FA_out_391+FA_cout_451;
  assign {FA_cout_1592,FA_out_1592}=FA_cout_391+FA_out_392+FA_cout_452;
  assign {FA_cout_1593,FA_out_1593}=FA_cout_392+FA_out_393+FA_cout_453;
  assign {FA_cout_1594,FA_out_1594}=FA_cout_393+FA_out_394+FA_cout_454;
  assign {FA_cout_1595,FA_out_1595}=FA_cout_394+FA_out_395+FA_cout_455;
  assign {FA_cout_1596,FA_out_1596}=FA_cout_395+FA_out_396+FA_cout_456;
  assign {FA_cout_1597,FA_out_1597}=FA_cout_396+FA_out_397+FA_cout_457;
  assign {FA_cout_1598,FA_out_1598}=FA_cout_397+FA_out_398+FA_cout_458;
  assign {FA_cout_1599,FA_out_1599}=FA_cout_398+FA_out_399+FA_cout_459;
  assign {FA_cout_1600,FA_out_1600}=FA_cout_399+FA_out_400+FA_cout_460;
  assign {FA_cout_1601,FA_out_1601}=FA_cout_400+FA_out_401+FA_cout_461;
  assign {FA_cout_1602,FA_out_1602}=FA_cout_401+FA_out_402+FA_cout_462;
  assign {FA_cout_1603,FA_out_1603}=FA_cout_402+FA_out_403+FA_cout_463;
  assign {FA_cout_1604,FA_out_1604}=FA_cout_403+FA_out_404+FA_cout_464;
  assign {FA_cout_1605,FA_out_1605}=FA_cout_404+FA_out_405+FA_cout_465;
  assign {FA_cout_1606,FA_out_1606}=FA_cout_405+FA_out_406+FA_cout_466;
  assign {FA_cout_1607,FA_out_1607}=FA_cout_406+FA_out_407+FA_cout_467;
  assign {FA_cout_1608,FA_out_1608}=FA_cout_407+FA_out_408+FA_cout_468;
  assign {FA_cout_1609,FA_out_1609}=FA_cout_408+FA_out_409+FA_cout_469;
  assign {FA_cout_1610,FA_out_1610}=FA_cout_409+FA_out_410+FA_cout_470;
  assign {FA_cout_1611,FA_out_1611}=FA_cout_410+FA_out_411+FA_cout_471;
  assign {FA_cout_1612,FA_out_1612}=FA_cout_411+FA_out_412+FA_cout_472;
  assign {FA_cout_1613,FA_out_1613}=FA_cout_412+FA_out_413+FA_cout_473;
  assign {FA_cout_1614,FA_out_1614}=FA_cout_413+FA_out_414+FA_cout_474;
  assign {FA_cout_1615,FA_out_1615}=FA_cout_414+FA_out_415+FA_cout_475;
  assign {FA_cout_1616,FA_out_1616}=FA_cout_415+FA_out_416+FA_cout_476;
  assign {FA_cout_1617,FA_out_1617}=FA_cout_416+FA_out_417+FA_cout_477;
  assign {FA_cout_1618,FA_out_1618}=FA_cout_417+FA_out_418+FA_cout_478;
  assign {FA_cout_1619,FA_out_1619}=FA_cout_418+FA_out_419+FA_cout_479;
  assign {FA_cout_1620,FA_out_1620}=FA_cout_419+FA_out_420+FA_cout_480;
  assign {FA_cout_1621,FA_out_1621}=FA_cout_420+FA_out_421+FA_cout_481;
  assign {FA_cout_1622,FA_out_1622}=FA_cout_421+FA_out_422+FA_cout_482;
  assign {FA_cout_1623,FA_out_1623}=FA_cout_422+FA_out_423+FA_cout_483;
  assign {FA_cout_1624,FA_out_1624}=FA_cout_423+FA_out_424+FA_cout_484;
  assign {FA_cout_1625,FA_out_1625}=FA_cout_424+FA_out_425+FA_cout_485;
  assign {FA_cout_1626,FA_out_1626}=FA_cout_425+FA_out_426+FA_cout_486;
  assign {FA_cout_1627,FA_out_1627}=FA_cout_426+FA_out_427+FA_cout_487;
  assign {FA_cout_1628,FA_out_1628}=FA_cout_427+FA_out_434+FA_cout_488;
  assign {FA_cout_1629,FA_out_1629}=FA_out_429+FA_cout_442+FA_out_490;
  assign {FA_cout_1630,FA_out_1630}=FA_cout_430+FA_out_437+FA_cout_491;
  assign {FA_cout_1631,FA_out_1631}=FA_out_432+FA_cout_445+FA_out_493;
  assign {FA_cout_1632,FA_out_1632}=FA_cout_433+FA_out_440+FA_cout_494;
  assign {FA_cout_1633,FA_out_1633}=FA_cout_434+FA_out_441+FA_cout_496;
  assign {FA_cout_1634,FA_out_1634}=FA_out_436+FA_cout_490+FA_out_498;
  assign {FA_cout_1635,FA_out_1635}=FA_cout_437+FA_out_444+FA_cout_499;
  assign {FA_cout_1636,FA_out_1636}=FA_out_439+FA_cout_493+FA_out_501;
  assign {FA_cout_1637,FA_out_1637}=FA_cout_440+FA_out_447+FA_cout_502;
  assign {FA_cout_1638,FA_out_1638}=FA_cout_441+FA_out_489+FA_cout_504;
  assign {FA_cout_1639,FA_out_1639}=FA_out_443+FA_cout_498+FA_out_506;
  assign {FA_cout_1640,FA_out_1640}=FA_cout_444+FA_out_492+FA_cout_507;
  assign {FA_cout_1641,FA_out_1641}=FA_out_446+FA_cout_501+FA_out_509;
  assign {FA_cout_1642,FA_out_1642}=FA_cout_447+FA_out_495+FA_cout_510;
  assign {FA_cout_1643,FA_out_1643}=FA_cout_489+FA_out_497+FA_cout_550;
  assign {FA_cout_1644,FA_out_1644}=FA_out_491+FA_cout_506+FA_out_552;
  assign {FA_cout_1645,FA_out_1645}=FA_cout_492+FA_out_500+FA_cout_553;
  assign {FA_cout_1646,FA_out_1646}=FA_out_494+FA_cout_509+FA_out_555;
  assign {FA_cout_1647,FA_out_1647}=FA_cout_495+FA_out_503+FA_cout_556;
  assign {FA_cout_1648,FA_out_1648}=FA_out_451+HA_cout_8+FA_out_512;
  assign {FA_cout_1649,FA_out_1649}=FA_out_452+FA_cout_512+FA_out_513;
  assign {FA_cout_1650,FA_out_1650}=FA_out_453+FA_cout_513+FA_out_514;
  assign {FA_cout_1651,FA_out_1651}=FA_out_454+FA_cout_514+FA_out_515;
  assign {FA_cout_1652,FA_out_1652}=FA_out_455+FA_cout_515+FA_out_516;
  assign {FA_cout_1653,FA_out_1653}=FA_out_456+FA_cout_516+FA_out_517;
  assign {FA_cout_1654,FA_out_1654}=FA_out_457+FA_cout_517+FA_out_518;
  assign {FA_cout_1655,FA_out_1655}=FA_out_458+FA_cout_518+FA_out_519;
  assign {FA_cout_1656,FA_out_1656}=FA_out_459+FA_cout_519+FA_out_520;
  assign {FA_cout_1657,FA_out_1657}=FA_out_460+FA_cout_520+FA_out_521;
  assign {FA_cout_1658,FA_out_1658}=FA_out_461+FA_cout_521+FA_out_522;
  assign {FA_cout_1659,FA_out_1659}=FA_out_462+FA_cout_522+FA_out_523;
  assign {FA_cout_1660,FA_out_1660}=FA_out_463+FA_cout_523+FA_out_524;
  assign {FA_cout_1661,FA_out_1661}=FA_out_464+FA_cout_524+FA_out_525;
  assign {FA_cout_1662,FA_out_1662}=FA_out_465+FA_cout_525+FA_out_526;
  assign {FA_cout_1663,FA_out_1663}=FA_out_466+FA_cout_526+FA_out_527;
  assign {FA_cout_1664,FA_out_1664}=FA_out_467+FA_cout_527+FA_out_528;
  assign {FA_cout_1665,FA_out_1665}=FA_out_468+FA_cout_528+FA_out_529;
  assign {FA_cout_1666,FA_out_1666}=FA_out_469+FA_cout_529+FA_out_530;
  assign {FA_cout_1667,FA_out_1667}=FA_out_470+FA_cout_530+FA_out_531;
  assign {FA_cout_1668,FA_out_1668}=FA_out_471+FA_cout_531+FA_out_532;
  assign {FA_cout_1669,FA_out_1669}=FA_out_472+FA_cout_532+FA_out_533;
  assign {FA_cout_1670,FA_out_1670}=FA_out_473+FA_cout_533+FA_out_534;
  assign {FA_cout_1671,FA_out_1671}=FA_out_474+FA_cout_534+FA_out_535;
  assign {FA_cout_1672,FA_out_1672}=FA_out_475+FA_cout_535+FA_out_536;
  assign {FA_cout_1673,FA_out_1673}=FA_out_476+FA_cout_536+FA_out_537;
  assign {FA_cout_1674,FA_out_1674}=FA_out_477+FA_cout_537+FA_out_538;
  assign {FA_cout_1675,FA_out_1675}=FA_out_478+FA_cout_538+FA_out_539;
  assign {FA_cout_1676,FA_out_1676}=FA_out_479+FA_cout_539+FA_out_540;
  assign {FA_cout_1677,FA_out_1677}=FA_out_480+FA_cout_540+FA_out_541;
  assign {FA_cout_1678,FA_out_1678}=FA_out_481+FA_cout_541+FA_out_542;
  assign {FA_cout_1679,FA_out_1679}=FA_out_482+FA_cout_542+FA_out_543;
  assign {FA_cout_1680,FA_out_1680}=FA_out_483+FA_cout_543+FA_out_544;
  assign {FA_cout_1681,FA_out_1681}=FA_out_484+FA_cout_544+FA_out_545;
  assign {FA_cout_1682,FA_out_1682}=FA_out_485+FA_cout_545+FA_out_546;
  assign {FA_cout_1683,FA_out_1683}=FA_out_486+FA_cout_546+FA_out_547;
  assign {FA_cout_1684,FA_out_1684}=FA_out_487+FA_cout_547+FA_out_548;
  assign {FA_cout_1685,FA_out_1685}=FA_out_488+FA_cout_548+FA_out_549;
  assign {FA_cout_1686,FA_out_1686}=FA_out_496+FA_cout_549+FA_out_558;
  assign {FA_cout_1687,FA_out_1687}=FA_cout_497+FA_out_505+FA_cout_559;
  assign {FA_cout_1688,FA_out_1688}=FA_out_499+FA_cout_552+FA_out_561;
  assign {FA_cout_1689,FA_out_1689}=FA_cout_500+FA_out_508+FA_cout_562;
  assign {FA_cout_1690,FA_out_1690}=FA_out_502+FA_cout_555+FA_out_564;
  assign {FA_cout_1691,FA_out_1691}=FA_cout_503+FA_out_511+FA_cout_565;
  assign {FA_cout_1692,FA_out_1692}=FA_out_504+FA_cout_558+FA_out_567;
  assign {FA_cout_1693,FA_out_1693}=FA_cout_505+FA_out_551+FA_cout_568;
  assign {FA_cout_1694,FA_out_1694}=FA_out_507+FA_cout_561+FA_out_570;
  assign {FA_cout_1695,FA_out_1695}=FA_cout_508+FA_out_554+FA_cout_571;
  assign {FA_cout_1696,FA_out_1696}=FA_out_510+FA_cout_564+FA_out_573;
  assign {FA_cout_1697,FA_out_1697}=FA_cout_511+FA_out_557+FA_cout_574;
  assign {FA_cout_1698,FA_out_1698}=FA_out_550+FA_cout_567+FA_out_611;
  assign {FA_cout_1699,FA_out_1699}=FA_cout_551+FA_out_560+FA_cout_612;
  assign {FA_cout_1700,FA_out_1700}=FA_out_553+FA_cout_570+FA_out_614;
  assign {FA_cout_1701,FA_out_1701}=FA_cout_554+FA_out_563+FA_cout_615;
  assign {FA_cout_1702,FA_out_1702}=FA_out_556+FA_cout_573+FA_out_617;
  assign {FA_cout_1703,FA_out_1703}=FA_cout_557+FA_out_566+FA_cout_618;
  assign {FA_cout_1704,FA_out_1704}=FA_out_559+FA_cout_611+FA_out_621;
  assign {FA_cout_1705,FA_out_1705}=FA_cout_560+FA_out_569+FA_cout_622;
  assign {FA_cout_1706,FA_out_1706}=FA_out_562+FA_cout_614+FA_out_624;
  assign {FA_cout_1707,FA_out_1707}=FA_cout_563+FA_out_572+FA_cout_625;
  assign {FA_cout_1708,FA_out_1708}=FA_out_565+FA_cout_617+FA_out_627;
  assign {FA_cout_1709,FA_out_1709}=FA_cout_566+FA_out_575+FA_cout_628;
  assign {FA_cout_1710,FA_out_1710}=FA_out_568+FA_cout_621+FA_out_631;
  assign {FA_cout_1711,FA_out_1711}=FA_cout_569+FA_out_613+FA_cout_632;
  assign {FA_cout_1712,FA_out_1712}=FA_out_571+FA_cout_624+FA_out_634;
  assign {FA_cout_1713,FA_out_1713}=FA_cout_572+FA_out_616+FA_cout_635;
  assign {FA_cout_1714,FA_out_1714}=FA_out_574+FA_cout_627+FA_out_637;
  assign {FA_cout_1715,FA_out_1715}=FA_cout_575+FA_out_619+FA_cout_638;
  assign {FA_cout_1716,FA_out_1716}=FA_cout_576+FA_out_577+inp_30[0];
  assign {FA_cout_1717,FA_out_1717}=FA_cout_577+FA_out_578+HA_out_10;
  assign {FA_cout_1718,FA_out_1718}=FA_cout_578+FA_out_579+HA_cout_10;
  assign {FA_cout_1719,FA_out_1719}=FA_cout_579+FA_out_580+FA_cout_640;
  assign {FA_cout_1720,FA_out_1720}=FA_cout_580+FA_out_581+FA_cout_641;
  assign {FA_cout_1721,FA_out_1721}=FA_cout_581+FA_out_582+FA_cout_642;
  assign {FA_cout_1722,FA_out_1722}=FA_cout_582+FA_out_583+FA_cout_643;
  assign {FA_cout_1723,FA_out_1723}=FA_cout_583+FA_out_584+FA_cout_644;
  assign {FA_cout_1724,FA_out_1724}=FA_cout_584+FA_out_585+FA_cout_645;
  assign {FA_cout_1725,FA_out_1725}=FA_cout_585+FA_out_586+FA_cout_646;
  assign {FA_cout_1726,FA_out_1726}=FA_cout_586+FA_out_587+FA_cout_647;
  assign {FA_cout_1727,FA_out_1727}=FA_cout_587+FA_out_588+FA_cout_648;
  assign {FA_cout_1728,FA_out_1728}=FA_cout_588+FA_out_589+FA_cout_649;
  assign {FA_cout_1729,FA_out_1729}=FA_cout_589+FA_out_590+FA_cout_650;
  assign {FA_cout_1730,FA_out_1730}=FA_cout_590+FA_out_591+FA_cout_651;
  assign {FA_cout_1731,FA_out_1731}=FA_cout_591+FA_out_592+FA_cout_652;
  assign {FA_cout_1732,FA_out_1732}=FA_cout_592+FA_out_593+FA_cout_653;
  assign {FA_cout_1733,FA_out_1733}=FA_cout_593+FA_out_594+FA_cout_654;
  assign {FA_cout_1734,FA_out_1734}=FA_cout_594+FA_out_595+FA_cout_655;
  assign {FA_cout_1735,FA_out_1735}=FA_cout_595+FA_out_596+FA_cout_656;
  assign {FA_cout_1736,FA_out_1736}=FA_cout_596+FA_out_597+FA_cout_657;
  assign {FA_cout_1737,FA_out_1737}=FA_cout_597+FA_out_598+FA_cout_658;
  assign {FA_cout_1738,FA_out_1738}=FA_cout_598+FA_out_599+FA_cout_659;
  assign {FA_cout_1739,FA_out_1739}=FA_cout_599+FA_out_600+FA_cout_660;
  assign {FA_cout_1740,FA_out_1740}=FA_cout_600+FA_out_601+FA_cout_661;
  assign {FA_cout_1741,FA_out_1741}=FA_cout_601+FA_out_602+FA_cout_662;
  assign {FA_cout_1742,FA_out_1742}=FA_cout_602+FA_out_603+FA_cout_663;
  assign {FA_cout_1743,FA_out_1743}=FA_cout_603+FA_out_604+FA_cout_664;
  assign {FA_cout_1744,FA_out_1744}=FA_cout_604+FA_out_605+FA_cout_665;
  assign {FA_cout_1745,FA_out_1745}=FA_cout_605+FA_out_606+FA_cout_666;
  assign {FA_cout_1746,FA_out_1746}=FA_cout_606+FA_out_607+FA_cout_667;
  assign {FA_cout_1747,FA_out_1747}=FA_cout_607+FA_out_608+FA_cout_668;
  assign {FA_cout_1748,FA_out_1748}=FA_cout_608+FA_out_609+FA_cout_669;
  assign {FA_cout_1749,FA_out_1749}=FA_cout_609+FA_out_610+FA_cout_670;
  assign {FA_cout_1750,FA_out_1750}=FA_cout_610+FA_out_620+FA_cout_671;
  assign {FA_cout_1751,FA_out_1751}=FA_out_612+FA_cout_631+FA_out_673;
  assign {FA_cout_1752,FA_out_1752}=FA_cout_613+FA_out_623+FA_cout_674;
  assign {FA_cout_1753,FA_out_1753}=FA_out_615+FA_cout_634+FA_out_676;
  assign {FA_cout_1754,FA_out_1754}=FA_cout_616+FA_out_626+FA_cout_677;
  assign {FA_cout_1755,FA_out_1755}=FA_out_618+FA_cout_637+FA_out_679;
  assign {FA_cout_1756,FA_out_1756}=FA_cout_619+FA_out_629+FA_cout_680;
  assign {FA_cout_1757,FA_out_1757}=FA_cout_620+FA_out_630+FA_cout_682;
  assign {FA_cout_1758,FA_out_1758}=FA_out_622+FA_cout_673+FA_out_684;
  assign {FA_cout_1759,FA_out_1759}=FA_cout_623+FA_out_633+FA_cout_685;
  assign {FA_cout_1760,FA_out_1760}=FA_out_625+FA_cout_676+FA_out_687;
  assign {FA_cout_1761,FA_out_1761}=FA_cout_626+FA_out_636+FA_cout_688;
  assign {FA_cout_1762,FA_out_1762}=FA_out_628+FA_cout_679+FA_out_690;
  assign {FA_cout_1763,FA_out_1763}=FA_cout_629+FA_out_639+FA_cout_691;
  assign {FA_cout_1764,FA_out_1764}=FA_cout_630+FA_out_672+FA_cout_693;
  assign {FA_cout_1765,FA_out_1765}=FA_out_632+FA_cout_684+FA_out_695;
  assign {FA_cout_1766,FA_out_1766}=FA_cout_633+FA_out_675+FA_cout_696;
  assign {FA_cout_1767,FA_out_1767}=FA_out_635+FA_cout_687+FA_out_698;
  assign {FA_cout_1768,FA_out_1768}=FA_cout_636+FA_out_678+FA_cout_699;
  assign {FA_cout_1769,FA_out_1769}=FA_out_638+FA_cout_690+FA_out_701;
  assign {FA_cout_1770,FA_out_1770}=FA_cout_639+FA_out_681+FA_cout_702;
  assign {FA_cout_1771,FA_out_1771}=FA_cout_672+FA_out_683+FA_cout_733;
  assign {FA_cout_1772,FA_out_1772}=FA_out_674+FA_cout_695+FA_out_735;
  assign {FA_cout_1773,FA_out_1773}=FA_cout_675+FA_out_686+FA_cout_736;
  assign {FA_cout_1774,FA_out_1774}=FA_out_677+FA_cout_698+FA_out_738;
  assign {FA_cout_1775,FA_out_1775}=FA_cout_678+FA_out_689+FA_cout_739;
  assign {FA_cout_1776,FA_out_1776}=FA_out_680+FA_cout_701+FA_out_741;
  assign {FA_cout_1777,FA_out_1777}=FA_cout_681+FA_out_692+FA_cout_742;
  assign {FA_cout_1778,FA_out_1778}=FA_out_643+HA_cout_11+FA_out_704;
  assign {FA_cout_1779,FA_out_1779}=FA_out_644+FA_cout_704+FA_out_705;
  assign {FA_cout_1780,FA_out_1780}=FA_out_645+FA_cout_705+FA_out_706;
  assign {FA_cout_1781,FA_out_1781}=FA_out_646+FA_cout_706+FA_out_707;
  assign {FA_cout_1782,FA_out_1782}=FA_out_647+FA_cout_707+FA_out_708;
  assign {FA_cout_1783,FA_out_1783}=FA_out_648+FA_cout_708+FA_out_709;
  assign {FA_cout_1784,FA_out_1784}=FA_out_649+FA_cout_709+FA_out_710;
  assign {FA_cout_1785,FA_out_1785}=FA_out_650+FA_cout_710+FA_out_711;
  assign {FA_cout_1786,FA_out_1786}=FA_out_651+FA_cout_711+FA_out_712;
  assign {FA_cout_1787,FA_out_1787}=FA_out_652+FA_cout_712+FA_out_713;
  assign {FA_cout_1788,FA_out_1788}=FA_out_653+FA_cout_713+FA_out_714;
  assign {FA_cout_1789,FA_out_1789}=FA_out_654+FA_cout_714+FA_out_715;
  assign {FA_cout_1790,FA_out_1790}=FA_out_655+FA_cout_715+FA_out_716;
  assign {FA_cout_1791,FA_out_1791}=FA_out_656+FA_cout_716+FA_out_717;
  assign {FA_cout_1792,FA_out_1792}=FA_out_657+FA_cout_717+FA_out_718;
  assign {FA_cout_1793,FA_out_1793}=FA_out_658+FA_cout_718+FA_out_719;
  assign {FA_cout_1794,FA_out_1794}=FA_out_659+FA_cout_719+FA_out_720;
  assign {FA_cout_1795,FA_out_1795}=FA_out_660+FA_cout_720+FA_out_721;
  assign {FA_cout_1796,FA_out_1796}=FA_out_661+FA_cout_721+FA_out_722;
  assign {FA_cout_1797,FA_out_1797}=FA_out_662+FA_cout_722+FA_out_723;
  assign {FA_cout_1798,FA_out_1798}=FA_out_663+FA_cout_723+FA_out_724;
  assign {FA_cout_1799,FA_out_1799}=FA_out_664+FA_cout_724+FA_out_725;
  assign {FA_cout_1800,FA_out_1800}=FA_out_665+FA_cout_725+FA_out_726;
  assign {FA_cout_1801,FA_out_1801}=FA_out_666+FA_cout_726+FA_out_727;
  assign {FA_cout_1802,FA_out_1802}=FA_out_667+FA_cout_727+FA_out_728;
  assign {FA_cout_1803,FA_out_1803}=FA_out_668+FA_cout_728+FA_out_729;
  assign {FA_cout_1804,FA_out_1804}=FA_out_669+FA_cout_729+FA_out_730;
  assign {FA_cout_1805,FA_out_1805}=FA_out_670+FA_cout_730+FA_out_731;
  assign {FA_cout_1806,FA_out_1806}=FA_out_671+FA_cout_731+FA_out_732;
  assign {FA_cout_1807,FA_out_1807}=FA_out_682+FA_cout_732+FA_out_744;
  assign {FA_cout_1808,FA_out_1808}=FA_cout_683+FA_out_694+FA_cout_745;
  assign {FA_cout_1809,FA_out_1809}=FA_out_685+FA_cout_735+FA_out_747;
  assign {FA_cout_1810,FA_out_1810}=FA_cout_686+FA_out_697+FA_cout_748;
  assign {FA_cout_1811,FA_out_1811}=FA_out_688+FA_cout_738+FA_out_750;
  assign {FA_cout_1812,FA_out_1812}=FA_cout_689+FA_out_700+FA_cout_751;
  assign {FA_cout_1813,FA_out_1813}=FA_out_691+FA_cout_741+FA_out_753;
  assign {FA_cout_1814,FA_out_1814}=FA_cout_692+FA_out_703+FA_cout_754;
  assign {FA_cout_1815,FA_out_1815}=FA_out_693+FA_cout_744+FA_out_756;
  assign {FA_cout_1816,FA_out_1816}=FA_cout_694+FA_out_734+FA_cout_757;
  assign {FA_cout_1817,FA_out_1817}=FA_out_696+FA_cout_747+FA_out_759;
  assign {FA_cout_1818,FA_out_1818}=FA_cout_697+FA_out_737+FA_cout_760;
  assign {FA_cout_1819,FA_out_1819}=FA_out_699+FA_cout_750+FA_out_762;
  assign {FA_cout_1820,FA_out_1820}=FA_cout_700+FA_out_740+FA_cout_763;
  assign {FA_cout_1821,FA_out_1821}=FA_out_702+FA_cout_753+FA_out_765;
  assign {FA_cout_1822,FA_out_1822}=FA_cout_703+FA_out_743+FA_cout_766;
  assign {FA_cout_1823,FA_out_1823}=FA_out_733+FA_cout_756+FA_out_794;
  assign {FA_cout_1824,FA_out_1824}=FA_cout_734+FA_out_746+FA_cout_795;
  assign {FA_cout_1825,FA_out_1825}=FA_out_736+FA_cout_759+FA_out_797;
  assign {FA_cout_1826,FA_out_1826}=FA_cout_737+FA_out_749+FA_cout_798;
  assign {FA_cout_1827,FA_out_1827}=FA_out_739+FA_cout_762+FA_out_800;
  assign {FA_cout_1828,FA_out_1828}=FA_cout_740+FA_out_752+FA_cout_801;
  assign {FA_cout_1829,FA_out_1829}=FA_out_742+FA_cout_765+FA_out_803;
  assign {FA_cout_1830,FA_out_1830}=FA_cout_743+FA_out_755+FA_cout_804;
  assign {FA_cout_1831,FA_out_1831}=FA_out_745+FA_cout_794+FA_out_807;
  assign {FA_cout_1832,FA_out_1832}=FA_cout_746+FA_out_758+FA_cout_808;
  assign {FA_cout_1833,FA_out_1833}=FA_out_748+FA_cout_797+FA_out_810;
  assign {FA_cout_1834,FA_out_1834}=FA_cout_749+FA_out_761+FA_cout_811;
  assign {FA_cout_1835,FA_out_1835}=FA_out_751+FA_cout_800+FA_out_813;
  assign {FA_cout_1836,FA_out_1836}=FA_cout_752+FA_out_764+FA_cout_814;
  assign {FA_cout_1837,FA_out_1837}=FA_out_754+FA_cout_803+FA_out_816;
  assign {FA_cout_1838,FA_out_1838}=FA_cout_755+FA_out_767+FA_cout_817;
  assign {FA_cout_1839,FA_out_1839}=FA_out_757+FA_cout_807+FA_out_820;
  assign {FA_cout_1840,FA_out_1840}=FA_cout_758+FA_out_796+FA_cout_821;
  assign {FA_cout_1841,FA_out_1841}=FA_out_760+FA_cout_810+FA_out_823;
  assign {FA_cout_1842,FA_out_1842}=FA_cout_761+FA_out_799+FA_cout_824;
  assign {FA_cout_1843,FA_out_1843}=FA_out_763+FA_cout_813+FA_out_826;
  assign {FA_cout_1844,FA_out_1844}=FA_cout_764+FA_out_802+FA_cout_827;
  assign {FA_cout_1845,FA_out_1845}=FA_out_766+FA_cout_816+FA_out_829;
  assign {FA_cout_1846,FA_out_1846}=FA_cout_767+FA_out_805+FA_cout_830;
  assign {FA_cout_1847,FA_out_1847}=FA_cout_768+FA_out_769+inp_39[0];
  assign {FA_cout_1848,FA_out_1848}=FA_cout_769+FA_out_770+HA_out_13;
  assign {FA_cout_1849,FA_out_1849}=FA_cout_770+FA_out_771+HA_cout_13;
  assign {FA_cout_1850,FA_out_1850}=FA_cout_771+FA_out_772+FA_cout_832;
  assign {FA_cout_1851,FA_out_1851}=FA_cout_772+FA_out_773+FA_cout_833;
  assign {FA_cout_1852,FA_out_1852}=FA_cout_773+FA_out_774+FA_cout_834;
  assign {FA_cout_1853,FA_out_1853}=FA_cout_774+FA_out_775+FA_cout_835;
  assign {FA_cout_1854,FA_out_1854}=FA_cout_775+FA_out_776+FA_cout_836;
  assign {FA_cout_1855,FA_out_1855}=FA_cout_776+FA_out_777+FA_cout_837;
  assign {FA_cout_1856,FA_out_1856}=FA_cout_777+FA_out_778+FA_cout_838;
  assign {FA_cout_1857,FA_out_1857}=FA_cout_778+FA_out_779+FA_cout_839;
  assign {FA_cout_1858,FA_out_1858}=FA_cout_779+FA_out_780+FA_cout_840;
  assign {FA_cout_1859,FA_out_1859}=FA_cout_780+FA_out_781+FA_cout_841;
  assign {FA_cout_1860,FA_out_1860}=FA_cout_781+FA_out_782+FA_cout_842;
  assign {FA_cout_1861,FA_out_1861}=FA_cout_782+FA_out_783+FA_cout_843;
  assign {FA_cout_1862,FA_out_1862}=FA_cout_783+FA_out_784+FA_cout_844;
  assign {FA_cout_1863,FA_out_1863}=FA_cout_784+FA_out_785+FA_cout_845;
  assign {FA_cout_1864,FA_out_1864}=FA_cout_785+FA_out_786+FA_cout_846;
  assign {FA_cout_1865,FA_out_1865}=FA_cout_786+FA_out_787+FA_cout_847;
  assign {FA_cout_1866,FA_out_1866}=FA_cout_787+FA_out_788+FA_cout_848;
  assign {FA_cout_1867,FA_out_1867}=FA_cout_788+FA_out_789+FA_cout_849;
  assign {FA_cout_1868,FA_out_1868}=FA_cout_789+FA_out_790+FA_cout_850;
  assign {FA_cout_1869,FA_out_1869}=FA_cout_790+FA_out_791+FA_cout_851;
  assign {FA_cout_1870,FA_out_1870}=FA_cout_791+FA_out_792+FA_cout_852;
  assign {FA_cout_1871,FA_out_1871}=FA_cout_792+FA_out_793+FA_cout_853;
  assign {FA_cout_1872,FA_out_1872}=FA_cout_793+FA_out_806+FA_cout_854;
  assign {FA_cout_1873,FA_out_1873}=FA_out_795+FA_cout_820+FA_out_856;
  assign {FA_cout_1874,FA_out_1874}=FA_cout_796+FA_out_809+FA_cout_857;
  assign {FA_cout_1875,FA_out_1875}=FA_out_798+FA_cout_823+FA_out_859;
  assign {FA_cout_1876,FA_out_1876}=FA_cout_799+FA_out_812+FA_cout_860;
  assign {FA_cout_1877,FA_out_1877}=FA_out_801+FA_cout_826+FA_out_862;
  assign {FA_cout_1878,FA_out_1878}=FA_cout_802+FA_out_815+FA_cout_863;
  assign {FA_cout_1879,FA_out_1879}=FA_out_804+FA_cout_829+FA_out_865;
  assign {FA_cout_1880,FA_out_1880}=FA_cout_805+FA_out_818+FA_cout_866;
  assign {FA_cout_1881,FA_out_1881}=FA_cout_806+FA_out_819+FA_cout_868;
  assign {FA_cout_1882,FA_out_1882}=FA_out_808+FA_cout_856+FA_out_870;
  assign {FA_cout_1883,FA_out_1883}=FA_cout_809+FA_out_822+FA_cout_871;
  assign {FA_cout_1884,FA_out_1884}=FA_out_811+FA_cout_859+FA_out_873;
  assign {FA_cout_1885,FA_out_1885}=FA_cout_812+FA_out_825+FA_cout_874;
  assign {FA_cout_1886,FA_out_1886}=FA_out_814+FA_cout_862+FA_out_876;
  assign {FA_cout_1887,FA_out_1887}=FA_cout_815+FA_out_828+FA_cout_877;
  assign {FA_cout_1888,FA_out_1888}=FA_out_817+FA_cout_865+FA_out_879;
  assign {FA_cout_1889,FA_out_1889}=FA_cout_818+FA_out_831+FA_cout_880;
  assign {FA_cout_1890,FA_out_1890}=FA_cout_819+FA_out_855+FA_cout_882;
  assign {FA_cout_1891,FA_out_1891}=FA_out_821+FA_cout_870+FA_out_884;
  assign {FA_cout_1892,FA_out_1892}=FA_cout_822+FA_out_858+FA_cout_885;
  assign {FA_cout_1893,FA_out_1893}=FA_out_824+FA_cout_873+FA_out_887;
  assign {FA_cout_1894,FA_out_1894}=FA_cout_825+FA_out_861+FA_cout_888;
  assign {FA_cout_1895,FA_out_1895}=FA_out_827+FA_cout_876+FA_out_890;
  assign {FA_cout_1896,FA_out_1896}=FA_cout_828+FA_out_864+FA_cout_891;
  assign {FA_cout_1897,FA_out_1897}=FA_out_830+FA_cout_879+FA_out_893;
  assign {FA_cout_1898,FA_out_1898}=FA_cout_831+FA_out_867+FA_cout_894;
  assign {FA_cout_1899,FA_out_1899}=FA_cout_855+FA_out_869+FA_cout_916;
  assign {FA_cout_1900,FA_out_1900}=FA_out_857+FA_cout_884+FA_out_918;
  assign {FA_cout_1901,FA_out_1901}=FA_cout_858+FA_out_872+FA_cout_919;
  assign {FA_cout_1902,FA_out_1902}=FA_out_860+FA_cout_887+FA_out_921;
  assign {FA_cout_1903,FA_out_1903}=FA_cout_861+FA_out_875+FA_cout_922;
  assign {FA_cout_1904,FA_out_1904}=FA_out_863+FA_cout_890+FA_out_924;
  assign {FA_cout_1905,FA_out_1905}=FA_cout_864+FA_out_878+FA_cout_925;
  assign {FA_cout_1906,FA_out_1906}=FA_out_866+FA_cout_893+FA_out_927;
  assign {FA_cout_1907,FA_out_1907}=FA_cout_867+FA_out_881+FA_cout_928;
  assign {FA_cout_1908,FA_out_1908}=FA_out_835+HA_cout_14+FA_out_896;
  assign {FA_cout_1909,FA_out_1909}=FA_out_836+FA_cout_896+FA_out_897;
  assign {FA_cout_1910,FA_out_1910}=FA_out_837+FA_cout_897+FA_out_898;
  assign {FA_cout_1911,FA_out_1911}=FA_out_838+FA_cout_898+FA_out_899;
  assign {FA_cout_1912,FA_out_1912}=FA_out_839+FA_cout_899+FA_out_900;
  assign {FA_cout_1913,FA_out_1913}=FA_out_840+FA_cout_900+FA_out_901;
  assign {FA_cout_1914,FA_out_1914}=FA_out_841+FA_cout_901+FA_out_902;
  assign {FA_cout_1915,FA_out_1915}=FA_out_842+FA_cout_902+FA_out_903;
  assign {FA_cout_1916,FA_out_1916}=FA_out_843+FA_cout_903+FA_out_904;
  assign {FA_cout_1917,FA_out_1917}=FA_out_844+FA_cout_904+FA_out_905;
  assign {FA_cout_1918,FA_out_1918}=FA_out_845+FA_cout_905+FA_out_906;
  assign {FA_cout_1919,FA_out_1919}=FA_out_846+FA_cout_906+FA_out_907;
  assign {FA_cout_1920,FA_out_1920}=FA_out_847+FA_cout_907+FA_out_908;
  assign {FA_cout_1921,FA_out_1921}=FA_out_848+FA_cout_908+FA_out_909;
  assign {FA_cout_1922,FA_out_1922}=FA_out_849+FA_cout_909+FA_out_910;
  assign {FA_cout_1923,FA_out_1923}=FA_out_850+FA_cout_910+FA_out_911;
  assign {FA_cout_1924,FA_out_1924}=FA_out_851+FA_cout_911+FA_out_912;
  assign {FA_cout_1925,FA_out_1925}=FA_out_852+FA_cout_912+FA_out_913;
  assign {FA_cout_1926,FA_out_1926}=FA_out_853+FA_cout_913+FA_out_914;
  assign {FA_cout_1927,FA_out_1927}=FA_out_854+FA_cout_914+FA_out_915;
  assign {FA_cout_1928,FA_out_1928}=FA_out_868+FA_cout_915+FA_out_930;
  assign {FA_cout_1929,FA_out_1929}=FA_cout_869+FA_out_883+FA_cout_931;
  assign {FA_cout_1930,FA_out_1930}=FA_out_871+FA_cout_918+FA_out_933;
  assign {FA_cout_1931,FA_out_1931}=FA_cout_872+FA_out_886+FA_cout_934;
  assign {FA_cout_1932,FA_out_1932}=FA_out_874+FA_cout_921+FA_out_936;
  assign {FA_cout_1933,FA_out_1933}=FA_cout_875+FA_out_889+FA_cout_937;
  assign {FA_cout_1934,FA_out_1934}=FA_out_877+FA_cout_924+FA_out_939;
  assign {FA_cout_1935,FA_out_1935}=FA_cout_878+FA_out_892+FA_cout_940;
  assign {FA_cout_1936,FA_out_1936}=FA_out_880+FA_cout_927+FA_out_942;
  assign {FA_cout_1937,FA_out_1937}=FA_cout_881+FA_out_895+FA_cout_943;
  assign {FA_cout_1938,FA_out_1938}=FA_out_882+FA_cout_930+FA_out_945;
  assign {FA_cout_1939,FA_out_1939}=FA_cout_883+FA_out_917+FA_cout_946;
  assign {FA_cout_1940,FA_out_1940}=FA_out_885+FA_cout_933+FA_out_948;
  assign {FA_cout_1941,FA_out_1941}=FA_cout_886+FA_out_920+FA_cout_949;
  assign {FA_cout_1942,FA_out_1942}=FA_out_888+FA_cout_936+FA_out_951;
  assign {FA_cout_1943,FA_out_1943}=FA_cout_889+FA_out_923+FA_cout_952;
  assign {FA_cout_1944,FA_out_1944}=FA_out_891+FA_cout_939+FA_out_954;
  assign {FA_cout_1945,FA_out_1945}=FA_cout_892+FA_out_926+FA_cout_955;
  assign {FA_cout_1946,FA_out_1946}=FA_out_894+FA_cout_942+FA_out_957;
  assign {FA_cout_1947,FA_out_1947}=FA_cout_895+FA_out_929+FA_cout_958;
  assign {FA_cout_1948,FA_out_1948}=FA_out_916+FA_cout_945+FA_out_977;
  assign {FA_cout_1949,FA_out_1949}=FA_cout_917+FA_out_932+FA_cout_978;
  assign {FA_cout_1950,FA_out_1950}=FA_out_919+FA_cout_948+FA_out_980;
  assign {FA_cout_1951,FA_out_1951}=FA_cout_920+FA_out_935+FA_cout_981;
  assign {FA_cout_1952,FA_out_1952}=FA_out_922+FA_cout_951+FA_out_983;
  assign {FA_cout_1953,FA_out_1953}=FA_cout_923+FA_out_938+FA_cout_984;
  assign {FA_cout_1954,FA_out_1954}=FA_out_925+FA_cout_954+FA_out_986;
  assign {FA_cout_1955,FA_out_1955}=FA_cout_926+FA_out_941+FA_cout_987;
  assign {FA_cout_1956,FA_out_1956}=FA_out_928+FA_cout_957+FA_out_989;
  assign {FA_cout_1957,FA_out_1957}=FA_cout_929+FA_out_944+FA_cout_990;
  assign {FA_cout_1958,FA_out_1958}=FA_out_931+FA_cout_977+FA_out_993;
  assign {FA_cout_1959,FA_out_1959}=FA_cout_932+FA_out_947+FA_cout_994;
  assign {FA_cout_1960,FA_out_1960}=FA_out_934+FA_cout_980+FA_out_996;
  assign {FA_cout_1961,FA_out_1961}=FA_cout_935+FA_out_950+FA_cout_997;
  assign {FA_cout_1962,FA_out_1962}=FA_out_937+FA_cout_983+FA_out_999;
  assign {FA_cout_1963,FA_out_1963}=FA_cout_938+FA_out_953+FA_cout_1000;
  assign {FA_cout_1964,FA_out_1964}=FA_out_940+FA_cout_986+FA_out_1002;
  assign {FA_cout_1965,FA_out_1965}=FA_cout_941+FA_out_956+FA_cout_1003;
  assign {FA_cout_1966,FA_out_1966}=FA_out_943+FA_cout_989+FA_out_1005;
  assign {FA_cout_1967,FA_out_1967}=FA_cout_944+FA_out_959+FA_cout_1006;
  assign {FA_cout_1968,FA_out_1968}=FA_out_946+FA_cout_993+FA_out_1009;
  assign {FA_cout_1969,FA_out_1969}=FA_cout_947+FA_out_979+FA_cout_1010;
  assign {FA_cout_1970,FA_out_1970}=FA_out_949+FA_cout_996+FA_out_1012;
  assign {FA_cout_1971,FA_out_1971}=FA_cout_950+FA_out_982+FA_cout_1013;
  assign {FA_cout_1972,FA_out_1972}=FA_out_952+FA_cout_999+FA_out_1015;
  assign {FA_cout_1973,FA_out_1973}=FA_cout_953+FA_out_985+FA_cout_1016;
  assign {FA_cout_1974,FA_out_1974}=FA_out_955+FA_cout_1002+FA_out_1018;
  assign {FA_cout_1975,FA_out_1975}=FA_cout_956+FA_out_988+FA_cout_1019;
  assign {FA_cout_1976,FA_out_1976}=FA_out_958+FA_cout_1005+FA_out_1021;
  assign {FA_cout_1977,FA_out_1977}=FA_cout_959+FA_out_991+FA_cout_1022;
  assign {FA_cout_1978,FA_out_1978}=FA_cout_960+FA_out_961+inp_48[0];
  assign {FA_cout_1979,FA_out_1979}=FA_cout_961+FA_out_962+HA_out_16;
  assign {FA_cout_1980,FA_out_1980}=FA_cout_962+FA_out_963+HA_cout_16;
  assign {FA_cout_1981,FA_out_1981}=FA_cout_963+FA_out_964+FA_cout_1024;
  assign {FA_cout_1982,FA_out_1982}=FA_cout_964+FA_out_965+FA_cout_1025;
  assign {FA_cout_1983,FA_out_1983}=FA_cout_965+FA_out_966+FA_cout_1026;
  assign {FA_cout_1984,FA_out_1984}=FA_cout_966+FA_out_967+FA_cout_1027;
  assign {FA_cout_1985,FA_out_1985}=FA_cout_967+FA_out_968+FA_cout_1028;
  assign {FA_cout_1986,FA_out_1986}=FA_cout_968+FA_out_969+FA_cout_1029;
  assign {FA_cout_1987,FA_out_1987}=FA_cout_969+FA_out_970+FA_cout_1030;
  assign {FA_cout_1988,FA_out_1988}=FA_cout_970+FA_out_971+FA_cout_1031;
  assign {FA_cout_1989,FA_out_1989}=FA_cout_971+FA_out_972+FA_cout_1032;
  assign {FA_cout_1990,FA_out_1990}=FA_cout_972+FA_out_973+FA_cout_1033;
  assign {FA_cout_1991,FA_out_1991}=FA_cout_973+FA_out_974+FA_cout_1034;
  assign {FA_cout_1992,FA_out_1992}=FA_cout_974+FA_out_975+FA_cout_1035;
  assign {FA_cout_1993,FA_out_1993}=FA_cout_975+FA_out_976+FA_cout_1036;
  assign {FA_cout_1994,FA_out_1994}=FA_cout_976+FA_out_992+FA_cout_1037;
  assign {FA_cout_1995,FA_out_1995}=FA_out_978+FA_cout_1009+FA_out_1039;
  assign {FA_cout_1996,FA_out_1996}=FA_cout_979+FA_out_995+FA_cout_1040;
  assign {FA_cout_1997,FA_out_1997}=FA_out_981+FA_cout_1012+FA_out_1042;
  assign {FA_cout_1998,FA_out_1998}=FA_cout_982+FA_out_998+FA_cout_1043;
  assign {FA_cout_1999,FA_out_1999}=FA_out_984+FA_cout_1015+FA_out_1045;
  assign {FA_cout_2000,FA_out_2000}=FA_cout_985+FA_out_1001+FA_cout_1046;
  assign {FA_cout_2001,FA_out_2001}=FA_out_987+FA_cout_1018+FA_out_1048;
  assign {FA_cout_2002,FA_out_2002}=FA_cout_988+FA_out_1004+FA_cout_1049;
  assign {FA_cout_2003,FA_out_2003}=FA_out_990+FA_cout_1021+FA_out_1051;
  assign {FA_cout_2004,FA_out_2004}=FA_cout_991+FA_out_1007+FA_cout_1052;
  assign {FA_cout_2005,FA_out_2005}=FA_cout_992+FA_out_1008+FA_cout_1054;
  assign {FA_cout_2006,FA_out_2006}=FA_out_994+FA_cout_1039+FA_out_1056;
  assign {FA_cout_2007,FA_out_2007}=FA_cout_995+FA_out_1011+FA_cout_1057;
  assign {FA_cout_2008,FA_out_2008}=FA_out_997+FA_cout_1042+FA_out_1059;
  assign {FA_cout_2009,FA_out_2009}=FA_cout_998+FA_out_1014+FA_cout_1060;
  assign {FA_cout_2010,FA_out_2010}=FA_out_1000+FA_cout_1045+FA_out_1062;
  assign {FA_cout_2011,FA_out_2011}=FA_cout_1001+FA_out_1017+FA_cout_1063;
  assign {FA_cout_2012,FA_out_2012}=FA_out_1003+FA_cout_1048+FA_out_1065;
  assign {FA_cout_2013,FA_out_2013}=FA_cout_1004+FA_out_1020+FA_cout_1066;
  assign {FA_cout_2014,FA_out_2014}=FA_out_1006+FA_cout_1051+FA_out_1068;
  assign {FA_cout_2015,FA_out_2015}=FA_cout_1007+FA_out_1023+FA_cout_1069;
  assign {FA_cout_2016,FA_out_2016}=FA_cout_1008+FA_out_1038+FA_cout_1071;
  assign {FA_cout_2017,FA_out_2017}=FA_out_1010+FA_cout_1056+FA_out_1073;
  assign {FA_cout_2018,FA_out_2018}=FA_cout_1011+FA_out_1041+FA_cout_1074;
  assign {FA_cout_2019,FA_out_2019}=FA_out_1013+FA_cout_1059+FA_out_1076;
  assign {FA_cout_2020,FA_out_2020}=FA_cout_1014+FA_out_1044+FA_cout_1077;
  assign {FA_cout_2021,FA_out_2021}=FA_out_1016+FA_cout_1062+FA_out_1079;
  assign {FA_cout_2022,FA_out_2022}=FA_cout_1017+FA_out_1047+FA_cout_1080;
  assign {FA_cout_2023,FA_out_2023}=FA_out_1019+FA_cout_1065+FA_out_1082;
  assign {FA_cout_2024,FA_out_2024}=FA_cout_1020+FA_out_1050+FA_cout_1083;
  assign {FA_cout_2025,FA_out_2025}=FA_out_1022+FA_cout_1068+FA_out_1085;
  assign {FA_cout_2026,FA_out_2026}=FA_cout_1023+FA_out_1053+FA_cout_1086;
  assign {FA_cout_2027,FA_out_2027}=FA_cout_1038+FA_out_1055+FA_cout_1099;
  assign {FA_cout_2028,FA_out_2028}=FA_out_1040+FA_cout_1073+FA_out_1101;
  assign {FA_cout_2029,FA_out_2029}=FA_cout_1041+FA_out_1058+FA_cout_1102;
  assign {FA_cout_2030,FA_out_2030}=FA_out_1043+FA_cout_1076+FA_out_1104;
  assign {FA_cout_2031,FA_out_2031}=FA_cout_1044+FA_out_1061+FA_cout_1105;
  assign {FA_cout_2032,FA_out_2032}=FA_out_1046+FA_cout_1079+FA_out_1107;
  assign {FA_cout_2033,FA_out_2033}=FA_cout_1047+FA_out_1064+FA_cout_1108;
  assign {FA_cout_2034,FA_out_2034}=FA_out_1049+FA_cout_1082+FA_out_1110;
  assign {FA_cout_2035,FA_out_2035}=FA_cout_1050+FA_out_1067+FA_cout_1111;
  assign {FA_cout_2036,FA_out_2036}=FA_out_1052+FA_cout_1085+FA_out_1113;
  assign {FA_cout_2037,FA_out_2037}=FA_cout_1053+FA_out_1070+FA_cout_1114;
  assign {FA_cout_2038,FA_out_2038}=FA_out_1027+HA_cout_17+FA_out_1088;
  assign {FA_cout_2039,FA_out_2039}=FA_out_1028+FA_cout_1088+FA_out_1089;
  assign {FA_cout_2040,FA_out_2040}=FA_out_1029+FA_cout_1089+FA_out_1090;
  assign {FA_cout_2041,FA_out_2041}=FA_out_1030+FA_cout_1090+FA_out_1091;
  assign {FA_cout_2042,FA_out_2042}=FA_out_1031+FA_cout_1091+FA_out_1092;
  assign {FA_cout_2043,FA_out_2043}=FA_out_1032+FA_cout_1092+FA_out_1093;
  assign {FA_cout_2044,FA_out_2044}=FA_out_1033+FA_cout_1093+FA_out_1094;
  assign {FA_cout_2045,FA_out_2045}=FA_out_1034+FA_cout_1094+FA_out_1095;
  assign {FA_cout_2046,FA_out_2046}=FA_out_1035+FA_cout_1095+FA_out_1096;
  assign {FA_cout_2047,FA_out_2047}=FA_out_1036+FA_cout_1096+FA_out_1097;
  assign {FA_cout_2048,FA_out_2048}=FA_out_1037+FA_cout_1097+FA_out_1098;
  assign {FA_cout_2049,FA_out_2049}=FA_out_1054+FA_cout_1098+FA_out_1116;
  assign {FA_cout_2050,FA_out_2050}=FA_cout_1055+FA_out_1072+FA_cout_1117;
  assign {FA_cout_2051,FA_out_2051}=FA_out_1057+FA_cout_1101+FA_out_1119;
  assign {FA_cout_2052,FA_out_2052}=FA_cout_1058+FA_out_1075+FA_cout_1120;
  assign {FA_cout_2053,FA_out_2053}=FA_out_1060+FA_cout_1104+FA_out_1122;
  assign {FA_cout_2054,FA_out_2054}=FA_cout_1061+FA_out_1078+FA_cout_1123;
  assign {FA_cout_2055,FA_out_2055}=FA_out_1063+FA_cout_1107+FA_out_1125;
  assign {FA_cout_2056,FA_out_2056}=FA_cout_1064+FA_out_1081+FA_cout_1126;
  assign {FA_cout_2057,FA_out_2057}=FA_out_1066+FA_cout_1110+FA_out_1128;
  assign {FA_cout_2058,FA_out_2058}=FA_cout_1067+FA_out_1084+FA_cout_1129;
  assign {FA_cout_2059,FA_out_2059}=FA_out_1069+FA_cout_1113+FA_out_1131;
  assign {FA_cout_2060,FA_out_2060}=FA_cout_1070+FA_out_1087+FA_cout_1132;
  assign {FA_cout_2061,FA_out_2061}=FA_out_1071+FA_cout_1116+FA_out_1134;
  assign {FA_cout_2062,FA_out_2062}=FA_cout_1072+FA_out_1100+FA_cout_1135;
  assign {FA_cout_2063,FA_out_2063}=FA_out_1074+FA_cout_1119+FA_out_1137;
  assign {FA_cout_2064,FA_out_2064}=FA_cout_1075+FA_out_1103+FA_cout_1138;
  assign {FA_cout_2065,FA_out_2065}=FA_out_1077+FA_cout_1122+FA_out_1140;
  assign {FA_cout_2066,FA_out_2066}=FA_cout_1078+FA_out_1106+FA_cout_1141;
  assign {FA_cout_2067,FA_out_2067}=FA_out_1080+FA_cout_1125+FA_out_1143;
  assign {FA_cout_2068,FA_out_2068}=FA_cout_1081+FA_out_1109+FA_cout_1144;
  assign {FA_cout_2069,FA_out_2069}=FA_out_1083+FA_cout_1128+FA_out_1146;
  assign {FA_cout_2070,FA_out_2070}=FA_cout_1084+FA_out_1112+FA_cout_1147;
  assign {FA_cout_2071,FA_out_2071}=FA_out_1086+FA_cout_1131+FA_out_1149;
  assign {FA_cout_2072,FA_out_2072}=FA_cout_1087+FA_out_1115+FA_cout_1150;
  assign {FA_cout_2073,FA_out_2073}=FA_out_1099+FA_cout_1134+FA_out_1160;
  assign {FA_cout_2074,FA_out_2074}=FA_cout_1100+FA_out_1118+FA_cout_1161;
  assign {FA_cout_2075,FA_out_2075}=FA_out_1102+FA_cout_1137+FA_out_1163;
  assign {FA_cout_2076,FA_out_2076}=FA_cout_1103+FA_out_1121+FA_cout_1164;
  assign {FA_cout_2077,FA_out_2077}=FA_out_1105+FA_cout_1140+FA_out_1166;
  assign {FA_cout_2078,FA_out_2078}=FA_cout_1106+FA_out_1124+FA_cout_1167;
  assign {FA_cout_2079,FA_out_2079}=FA_out_1108+FA_cout_1143+FA_out_1169;
  assign {FA_cout_2080,FA_out_2080}=FA_cout_1109+FA_out_1127+FA_cout_1170;
  assign {FA_cout_2081,FA_out_2081}=FA_out_1111+FA_cout_1146+FA_out_1172;
  assign {FA_cout_2082,FA_out_2082}=FA_cout_1112+FA_out_1130+FA_cout_1173;
  assign {FA_cout_2083,FA_out_2083}=FA_out_1114+FA_cout_1149+FA_out_1175;
  assign {FA_cout_2084,FA_out_2084}=FA_cout_1115+FA_out_1133+FA_cout_1176;
  assign {FA_cout_2085,FA_out_2085}=FA_out_1117+FA_cout_1160+FA_out_1179;
  assign {FA_cout_2086,FA_out_2086}=FA_cout_1118+FA_out_1136+FA_cout_1180;
  assign {FA_cout_2087,FA_out_2087}=FA_out_1120+FA_cout_1163+FA_out_1182;
  assign {FA_cout_2088,FA_out_2088}=FA_cout_1121+FA_out_1139+FA_cout_1183;
  assign {FA_cout_2089,FA_out_2089}=FA_out_1123+FA_cout_1166+FA_out_1185;
  assign {FA_cout_2090,FA_out_2090}=FA_cout_1124+FA_out_1142+FA_cout_1186;
  assign {FA_cout_2091,FA_out_2091}=FA_out_1126+FA_cout_1169+FA_out_1188;
  assign {FA_cout_2092,FA_out_2092}=FA_cout_1127+FA_out_1145+FA_cout_1189;
  assign {FA_cout_2093,FA_out_2093}=FA_out_1129+FA_cout_1172+FA_out_1191;
  assign {FA_cout_2094,FA_out_2094}=FA_cout_1130+FA_out_1148+FA_cout_1192;
  assign {FA_cout_2095,FA_out_2095}=FA_out_1132+FA_cout_1175+FA_out_1194;
  assign {FA_cout_2096,FA_out_2096}=FA_cout_1133+FA_out_1151+FA_cout_1195;
  assign {FA_cout_2097,FA_out_2097}=FA_out_1135+FA_cout_1179+FA_out_1198;
  assign {FA_cout_2098,FA_out_2098}=FA_cout_1136+FA_out_1162+FA_cout_1199;
  assign {FA_cout_2099,FA_out_2099}=FA_out_1138+FA_cout_1182+FA_out_1201;
  assign {FA_cout_2100,FA_out_2100}=FA_cout_1139+FA_out_1165+FA_cout_1202;
  assign {FA_cout_2101,FA_out_2101}=FA_out_1141+FA_cout_1185+FA_out_1204;
  assign {FA_cout_2102,FA_out_2102}=FA_cout_1142+FA_out_1168+FA_cout_1205;
  assign {FA_cout_2103,FA_out_2103}=FA_out_1144+FA_cout_1188+FA_out_1207;
  assign {FA_cout_2104,FA_out_2104}=FA_cout_1145+FA_out_1171+FA_cout_1208;
  assign {FA_cout_2105,FA_out_2105}=FA_out_1147+FA_cout_1191+FA_out_1210;
  assign {FA_cout_2106,FA_out_2106}=FA_cout_1148+FA_out_1174+FA_cout_1211;
  assign {FA_cout_2107,FA_out_2107}=FA_out_1150+FA_cout_1194+FA_out_1213;
  assign {FA_cout_2108,FA_out_2108}=FA_cout_1151+FA_out_1177+FA_cout_1214;
  assign {FA_cout_2109,FA_out_2109}=FA_cout_1152+FA_out_1153+inp_57[0];
  assign {FA_cout_2110,FA_out_2110}=FA_cout_1153+FA_out_1154+HA_out_19;
  assign {FA_cout_2111,FA_out_2111}=FA_cout_1154+FA_out_1155+HA_cout_19;
  assign {FA_cout_2112,FA_out_2112}=FA_cout_1155+FA_out_1156+FA_cout_1216;
  assign {FA_cout_2113,FA_out_2113}=FA_cout_1156+FA_out_1157+FA_cout_1217;
  assign {FA_cout_2114,FA_out_2114}=FA_cout_1157+FA_out_1158+FA_cout_1218;
  assign {FA_cout_2115,FA_out_2115}=FA_cout_1158+FA_out_1159+FA_cout_1219;
  assign {FA_cout_2116,FA_out_2116}=FA_cout_1159+FA_out_1178+FA_cout_1220;
  assign {FA_cout_2117,FA_out_2117}=FA_out_1161+FA_cout_1198+FA_out_1222;
  assign {FA_cout_2118,FA_out_2118}=FA_cout_1162+FA_out_1181+FA_cout_1223;
  assign {FA_cout_2119,FA_out_2119}=FA_out_1164+FA_cout_1201+FA_out_1225;
  assign {FA_cout_2120,FA_out_2120}=FA_cout_1165+FA_out_1184+FA_cout_1226;
  assign {FA_cout_2121,FA_out_2121}=FA_out_1167+FA_cout_1204+FA_out_1228;
  assign {FA_cout_2122,FA_out_2122}=FA_cout_1168+FA_out_1187+FA_cout_1229;
  assign {FA_cout_2123,FA_out_2123}=FA_out_1170+FA_cout_1207+FA_out_1231;
  assign {FA_cout_2124,FA_out_2124}=FA_cout_1171+FA_out_1190+FA_cout_1232;
  assign {FA_cout_2125,FA_out_2125}=FA_out_1173+FA_cout_1210+FA_out_1234;
  assign {FA_cout_2126,FA_out_2126}=FA_cout_1174+FA_out_1193+FA_cout_1235;
  assign {FA_cout_2127,FA_out_2127}=FA_out_1176+FA_cout_1213+FA_out_1237;
  assign {FA_cout_2128,FA_out_2128}=FA_cout_1177+FA_out_1196+FA_cout_1238;
  assign {FA_cout_2129,FA_out_2129}=FA_cout_1178+FA_out_1197+FA_cout_1240;
  assign {FA_cout_2130,FA_out_2130}=FA_out_1180+FA_cout_1222+FA_out_1242;
  assign {FA_cout_2131,FA_out_2131}=FA_cout_1181+FA_out_1200+FA_cout_1243;
  assign {FA_cout_2132,FA_out_2132}=FA_out_1183+FA_cout_1225+FA_out_1245;
  assign {FA_cout_2133,FA_out_2133}=FA_cout_1184+FA_out_1203+FA_cout_1246;
  assign {FA_cout_2134,FA_out_2134}=FA_out_1186+FA_cout_1228+FA_out_1248;
  assign {FA_cout_2135,FA_out_2135}=FA_cout_1187+FA_out_1206+FA_cout_1249;
  assign {FA_cout_2136,FA_out_2136}=FA_out_1189+FA_cout_1231+FA_out_1251;
  assign {FA_cout_2137,FA_out_2137}=FA_cout_1190+FA_out_1209+FA_cout_1252;
  assign {FA_cout_2138,FA_out_2138}=FA_out_1192+FA_cout_1234+FA_out_1254;
  assign {FA_cout_2139,FA_out_2139}=FA_cout_1193+FA_out_1212+FA_cout_1255;
  assign {FA_cout_2140,FA_out_2140}=FA_out_1195+FA_cout_1237+FA_out_1257;
  assign {FA_cout_2141,FA_out_2141}=FA_cout_1196+FA_out_1215+FA_cout_1258;
  assign {FA_cout_2142,FA_out_2142}=FA_cout_1197+FA_out_1221+FA_cout_1260;
  assign {FA_cout_2143,FA_out_2143}=FA_out_1199+FA_cout_1242+FA_out_1262;
  assign {FA_cout_2144,FA_out_2144}=FA_cout_1200+FA_out_1224+FA_cout_1263;
  assign {FA_cout_2145,FA_out_2145}=FA_out_1202+FA_cout_1245+FA_out_1265;
  assign {FA_cout_2146,FA_out_2146}=FA_cout_1203+FA_out_1227+FA_cout_1266;
  assign {FA_cout_2147,FA_out_2147}=FA_out_1205+FA_cout_1248+FA_out_1268;
  assign {FA_cout_2148,FA_out_2148}=FA_cout_1206+FA_out_1230+FA_cout_1269;
  assign {FA_cout_2149,FA_out_2149}=FA_out_1208+FA_cout_1251+FA_out_1271;
  assign {FA_cout_2150,FA_out_2150}=FA_cout_1209+FA_out_1233+FA_cout_1272;
  assign {FA_cout_2151,FA_out_2151}=FA_out_1211+FA_cout_1254+FA_out_1274;
  assign {FA_cout_2152,FA_out_2152}=FA_cout_1212+FA_out_1236+FA_cout_1275;
  assign {FA_cout_2153,FA_out_2153}=FA_out_1214+FA_cout_1257+FA_out_1277;
  assign {FA_cout_2154,FA_out_2154}=FA_cout_1215+FA_out_1239+FA_cout_1278;
  assign {FA_cout_2155,FA_out_2155}=FA_cout_1221+FA_out_1241+FA_cout_1282;
  assign {FA_cout_2156,FA_out_2156}=FA_out_1223+FA_cout_1262+FA_out_1284;
  assign {FA_cout_2157,FA_out_2157}=FA_cout_1224+FA_out_1244+FA_cout_1285;
  assign {FA_cout_2158,FA_out_2158}=FA_out_1226+FA_cout_1265+FA_out_1287;
  assign {FA_cout_2159,FA_out_2159}=FA_cout_1227+FA_out_1247+FA_cout_1288;
  assign {FA_cout_2160,FA_out_2160}=FA_out_1229+FA_cout_1268+FA_out_1290;
  assign {FA_cout_2161,FA_out_2161}=FA_cout_1230+FA_out_1250+FA_cout_1291;
  assign {FA_cout_2162,FA_out_2162}=FA_out_1232+FA_cout_1271+FA_out_1293;
  assign {FA_cout_2163,FA_out_2163}=FA_cout_1233+FA_out_1253+FA_cout_1294;
  assign {FA_cout_2164,FA_out_2164}=FA_out_1235+FA_cout_1274+FA_out_1296;
  assign {FA_cout_2165,FA_out_2165}=FA_cout_1236+FA_out_1256+FA_cout_1297;
  assign {FA_cout_2166,FA_out_2166}=FA_out_1238+FA_cout_1277+FA_out_1299;
  assign {FA_cout_2167,FA_out_2167}=FA_cout_1239+FA_out_1259+FA_cout_1300;
  assign {FA_cout_2168,FA_out_2168}=FA_out_1219+HA_cout_20+FA_out_1280;
  assign {FA_cout_2169,FA_out_2169}=FA_out_1220+FA_cout_1280+FA_out_1281;
  assign {FA_cout_2170,FA_out_2170}=FA_out_1240+FA_cout_1281+FA_out_1302;
  assign {FA_cout_2171,FA_out_2171}=FA_cout_1241+FA_out_1261+FA_cout_1303;
  assign {FA_cout_2172,FA_out_2172}=FA_out_1243+FA_cout_1284+FA_out_1305;
  assign {FA_cout_2173,FA_out_2173}=FA_cout_1244+FA_out_1264+FA_cout_1306;
  assign {FA_cout_2174,FA_out_2174}=FA_out_1246+FA_cout_1287+FA_out_1308;
  assign {FA_cout_2175,FA_out_2175}=FA_cout_1247+FA_out_1267+FA_cout_1309;
  assign {FA_cout_2176,FA_out_2176}=FA_out_1249+FA_cout_1290+FA_out_1311;
  assign {FA_cout_2177,FA_out_2177}=FA_cout_1250+FA_out_1270+FA_cout_1312;
  assign {FA_cout_2178,FA_out_2178}=FA_out_1252+FA_cout_1293+FA_out_1314;
  assign {FA_cout_2179,FA_out_2179}=FA_cout_1253+FA_out_1273+FA_cout_1315;
  assign {FA_cout_2180,FA_out_2180}=FA_out_1255+FA_cout_1296+FA_out_1317;
  assign {FA_cout_2181,FA_out_2181}=FA_cout_1256+FA_out_1276+FA_cout_1318;
  assign {FA_cout_2182,FA_out_2182}=FA_out_1258+FA_cout_1299+FA_out_1320;
  assign {FA_cout_2183,FA_out_2183}=FA_cout_1259+FA_out_1279+FA_cout_1321;
  assign {FA_cout_2184,FA_out_2184}=FA_out_1260+FA_cout_1302+HA_out_21;
  assign {FA_cout_2185,FA_out_2185}=FA_cout_1261+FA_out_1283+HA_cout_22;
  assign {FA_cout_2186,FA_out_2186}=FA_out_1263+FA_cout_1305+HA_out_24;
  assign {FA_cout_2187,FA_out_2187}=FA_cout_1264+FA_out_1286+HA_cout_25;
  assign {FA_cout_2188,FA_out_2188}=FA_out_1266+FA_cout_1308+HA_out_27;
  assign {FA_cout_2189,FA_out_2189}=FA_cout_1267+FA_out_1289+HA_cout_28;
  assign {FA_cout_2190,FA_out_2190}=FA_out_1269+FA_cout_1311+HA_out_30;
  assign {FA_cout_2191,FA_out_2191}=FA_cout_1270+FA_out_1292+HA_cout_31;
  assign {FA_cout_2192,FA_out_2192}=FA_out_1272+FA_cout_1314+HA_out_33;
  assign {FA_cout_2193,FA_out_2193}=FA_cout_1273+FA_out_1295+HA_cout_34;
  assign {FA_cout_2194,FA_out_2194}=FA_out_1275+FA_cout_1317+HA_out_36;
  assign {FA_cout_2195,FA_out_2195}=FA_cout_1276+FA_out_1298+HA_cout_37;
  assign {FA_cout_2196,FA_out_2196}=FA_out_1278+FA_cout_1320+HA_out_39;
  assign {FA_cout_2197,FA_out_2197}=FA_cout_1279+FA_out_1301+HA_cout_40;
  assign {FA_cout_2198,FA_out_2198}=FA_out_1282+HA_cout_21+inp_63[3];
  assign {FA_cout_2199,FA_out_2199}=FA_out_1285+HA_cout_24+inp_63[12];
  assign {FA_cout_2200,FA_out_2200}=FA_out_1288+HA_cout_27+inp_63[21];
  assign {FA_cout_2201,FA_out_2201}=FA_out_1291+HA_cout_30+inp_63[30];
  assign {FA_cout_2202,FA_out_2202}=FA_out_1294+HA_cout_33+inp_63[39];
  assign {FA_cout_2203,FA_out_2203}=FA_out_1297+HA_cout_36+inp_63[48];
  assign {FA_cout_2204,FA_out_2204}=FA_out_1300+HA_cout_39+inp_63[57];
  assign {FA_cout_2205,FA_out_2205}=FA_cout_1324+FA_out_1325+FA_out_64;
  assign {FA_cout_2206,FA_out_2206}=FA_cout_1325+FA_out_1326+HA_out_43;
  assign {FA_cout_2207,FA_out_2207}=FA_cout_1326+FA_out_1327+HA_cout_43;
  assign {FA_cout_2208,FA_out_2208}=FA_cout_1327+FA_out_1328+HA_cout_44;
  assign {FA_cout_2209,FA_out_2209}=FA_cout_1328+FA_out_1329+FA_cout_1388;
  assign {FA_cout_2210,FA_out_2210}=FA_cout_1329+FA_out_1330+FA_cout_1389;
  assign {FA_cout_2211,FA_out_2211}=FA_cout_1330+FA_out_1331+FA_cout_1390;
  assign {FA_cout_2212,FA_out_2212}=FA_cout_1331+FA_out_1332+FA_cout_1391;
  assign {FA_cout_2213,FA_out_2213}=FA_cout_1332+FA_out_1333+FA_cout_1392;
  assign {FA_cout_2214,FA_out_2214}=FA_cout_1333+FA_out_1334+FA_cout_1393;
  assign {FA_cout_2215,FA_out_2215}=FA_cout_1334+FA_out_1335+FA_cout_1394;
  assign {FA_cout_2216,FA_out_2216}=FA_cout_1335+FA_out_1336+FA_cout_1395;
  assign {FA_cout_2217,FA_out_2217}=FA_cout_1336+FA_out_1337+FA_cout_1396;
  assign {FA_cout_2218,FA_out_2218}=FA_cout_1337+FA_out_1338+FA_cout_1397;
  assign {FA_cout_2219,FA_out_2219}=FA_cout_1338+FA_out_1339+FA_cout_1398;
  assign {FA_cout_2220,FA_out_2220}=FA_cout_1339+FA_out_1340+FA_cout_1399;
  assign {FA_cout_2221,FA_out_2221}=FA_cout_1340+FA_out_1341+FA_cout_1400;
  assign {FA_cout_2222,FA_out_2222}=FA_cout_1341+FA_out_1342+FA_cout_1401;
  assign {FA_cout_2223,FA_out_2223}=FA_cout_1342+FA_out_1343+FA_cout_1402;
  assign {FA_cout_2224,FA_out_2224}=FA_cout_1343+FA_out_1344+FA_cout_1403;
  assign {FA_cout_2225,FA_out_2225}=FA_cout_1344+FA_out_1345+FA_cout_1404;
  assign {FA_cout_2226,FA_out_2226}=FA_cout_1345+FA_out_1346+FA_cout_1405;
  assign {FA_cout_2227,FA_out_2227}=FA_cout_1346+FA_out_1347+FA_cout_1406;
  assign {FA_cout_2228,FA_out_2228}=FA_cout_1347+FA_out_1348+FA_cout_1407;
  assign {FA_cout_2229,FA_out_2229}=FA_cout_1348+FA_out_1349+FA_cout_1408;
  assign {FA_cout_2230,FA_out_2230}=FA_cout_1349+FA_out_1350+FA_cout_1409;
  assign {FA_cout_2231,FA_out_2231}=FA_cout_1350+FA_out_1351+FA_cout_1410;
  assign {FA_cout_2232,FA_out_2232}=FA_cout_1351+FA_out_1352+FA_cout_1411;
  assign {FA_cout_2233,FA_out_2233}=FA_cout_1352+FA_out_1353+FA_cout_1412;
  assign {FA_cout_2234,FA_out_2234}=FA_cout_1353+FA_out_1354+FA_cout_1413;
  assign {FA_cout_2235,FA_out_2235}=FA_cout_1354+FA_out_1355+FA_cout_1414;
  assign {FA_cout_2236,FA_out_2236}=FA_cout_1355+FA_out_1356+FA_cout_1415;
  assign {FA_cout_2237,FA_out_2237}=FA_cout_1356+FA_out_1357+FA_cout_1416;
  assign {FA_cout_2238,FA_out_2238}=FA_cout_1357+FA_out_1358+FA_cout_1417;
  assign {FA_cout_2239,FA_out_2239}=FA_cout_1358+FA_out_1359+FA_cout_1418;
  assign {FA_cout_2240,FA_out_2240}=FA_cout_1359+FA_out_1360+FA_cout_1419;
  assign {FA_cout_2241,FA_out_2241}=FA_cout_1360+FA_out_1361+FA_cout_1420;
  assign {FA_cout_2242,FA_out_2242}=FA_cout_1361+FA_out_1362+FA_cout_1421;
  assign {FA_cout_2243,FA_out_2243}=FA_cout_1362+FA_out_1363+FA_cout_1422;
  assign {FA_cout_2244,FA_out_2244}=FA_cout_1363+FA_out_1364+FA_cout_1423;
  assign {FA_cout_2245,FA_out_2245}=FA_cout_1364+FA_out_1365+FA_cout_1424;
  assign {FA_cout_2246,FA_out_2246}=FA_cout_1365+FA_out_1366+FA_cout_1425;
  assign {FA_cout_2247,FA_out_2247}=FA_cout_1366+FA_out_1367+FA_cout_1426;
  assign {FA_cout_2248,FA_out_2248}=FA_cout_1367+FA_out_1368+FA_cout_1427;
  assign {FA_cout_2249,FA_out_2249}=FA_cout_1368+FA_out_1369+FA_cout_1428;
  assign {FA_cout_2250,FA_out_2250}=FA_cout_1369+FA_out_1370+FA_cout_1429;
  assign {FA_cout_2251,FA_out_2251}=FA_cout_1370+FA_out_1371+FA_cout_1430;
  assign {FA_cout_2252,FA_out_2252}=FA_cout_1371+FA_out_1372+FA_cout_1431;
  assign {FA_cout_2253,FA_out_2253}=FA_cout_1372+FA_out_1373+FA_cout_1432;
  assign {FA_cout_2254,FA_out_2254}=FA_cout_1373+FA_out_1374+FA_cout_1433;
  assign {FA_cout_2255,FA_out_2255}=FA_cout_1374+FA_out_1375+FA_cout_1434;
  assign {FA_cout_2256,FA_out_2256}=FA_cout_1375+FA_out_1376+FA_cout_1435;
  assign {FA_cout_2257,FA_out_2257}=FA_cout_1376+FA_out_1377+FA_cout_1436;
  assign {FA_cout_2258,FA_out_2258}=FA_cout_1377+FA_out_1378+FA_cout_1437;
  assign {FA_cout_2259,FA_out_2259}=FA_cout_1378+FA_out_1379+FA_cout_1438;
  assign {FA_cout_2260,FA_out_2260}=FA_cout_1379+FA_out_1380+FA_cout_1439;
  assign {FA_cout_2261,FA_out_2261}=FA_cout_1380+FA_out_1381+FA_cout_1440;
  assign {FA_cout_2262,FA_out_2262}=FA_cout_1381+FA_out_1382+FA_cout_1441;
  assign {FA_cout_2263,FA_out_2263}=FA_cout_1382+FA_out_1383+FA_cout_1442;
  assign {FA_cout_2264,FA_out_2264}=FA_cout_1383+FA_out_1384+FA_cout_1443;
  assign {FA_cout_2265,FA_out_2265}=FA_cout_1384+FA_out_1385+FA_cout_1444;
  assign {FA_cout_2266,FA_out_2266}=FA_cout_1385+FA_out_1386+FA_cout_1446;
  assign {FA_cout_2267,FA_out_2267}=FA_cout_1386+FA_out_1387+FA_cout_1448;
  assign {FA_cout_2268,FA_out_2268}=FA_cout_1387+FA_out_1445+FA_cout_1450;
  assign {FA_cout_2269,FA_out_2269}=FA_cout_1445+FA_out_1447+FA_cout_1452;
  assign {FA_cout_2270,FA_out_2270}=FA_out_1392+HA_cout_45+FA_out_1454;
  assign {FA_cout_2271,FA_out_2271}=FA_out_1393+FA_cout_1454+FA_out_1455;
  assign {FA_cout_2272,FA_out_2272}=FA_out_1394+FA_cout_1455+FA_out_1456;
  assign {FA_cout_2273,FA_out_2273}=FA_out_1395+FA_cout_1456+FA_out_1457;
  assign {FA_cout_2274,FA_out_2274}=FA_out_1396+FA_cout_1457+FA_out_1458;
  assign {FA_cout_2275,FA_out_2275}=FA_out_1397+FA_cout_1458+FA_out_1459;
  assign {FA_cout_2276,FA_out_2276}=FA_out_1398+FA_cout_1459+FA_out_1460;
  assign {FA_cout_2277,FA_out_2277}=FA_out_1399+FA_cout_1460+FA_out_1461;
  assign {FA_cout_2278,FA_out_2278}=FA_out_1400+FA_cout_1461+FA_out_1462;
  assign {FA_cout_2279,FA_out_2279}=FA_out_1401+FA_cout_1462+FA_out_1463;
  assign {FA_cout_2280,FA_out_2280}=FA_out_1402+FA_cout_1463+FA_out_1464;
  assign {FA_cout_2281,FA_out_2281}=FA_out_1403+FA_cout_1464+FA_out_1465;
  assign {FA_cout_2282,FA_out_2282}=FA_out_1404+FA_cout_1465+FA_out_1466;
  assign {FA_cout_2283,FA_out_2283}=FA_out_1405+FA_cout_1466+FA_out_1467;
  assign {FA_cout_2284,FA_out_2284}=FA_out_1406+FA_cout_1467+FA_out_1468;
  assign {FA_cout_2285,FA_out_2285}=FA_out_1407+FA_cout_1468+FA_out_1469;
  assign {FA_cout_2286,FA_out_2286}=FA_out_1408+FA_cout_1469+FA_out_1470;
  assign {FA_cout_2287,FA_out_2287}=FA_out_1409+FA_cout_1470+FA_out_1471;
  assign {FA_cout_2288,FA_out_2288}=FA_out_1410+FA_cout_1471+FA_out_1472;
  assign {FA_cout_2289,FA_out_2289}=FA_out_1411+FA_cout_1472+FA_out_1473;
  assign {FA_cout_2290,FA_out_2290}=FA_out_1412+FA_cout_1473+FA_out_1474;
  assign {FA_cout_2291,FA_out_2291}=FA_out_1413+FA_cout_1474+FA_out_1475;
  assign {FA_cout_2292,FA_out_2292}=FA_out_1414+FA_cout_1475+FA_out_1476;
  assign {FA_cout_2293,FA_out_2293}=FA_out_1415+FA_cout_1476+FA_out_1477;
  assign {FA_cout_2294,FA_out_2294}=FA_out_1416+FA_cout_1477+FA_out_1478;
  assign {FA_cout_2295,FA_out_2295}=FA_out_1417+FA_cout_1478+FA_out_1479;
  assign {FA_cout_2296,FA_out_2296}=FA_out_1418+FA_cout_1479+FA_out_1480;
  assign {FA_cout_2297,FA_out_2297}=FA_out_1419+FA_cout_1480+FA_out_1481;
  assign {FA_cout_2298,FA_out_2298}=FA_out_1420+FA_cout_1481+FA_out_1482;
  assign {FA_cout_2299,FA_out_2299}=FA_out_1421+FA_cout_1482+FA_out_1483;
  assign {FA_cout_2300,FA_out_2300}=FA_out_1422+FA_cout_1483+FA_out_1484;
  assign {FA_cout_2301,FA_out_2301}=FA_out_1423+FA_cout_1484+FA_out_1485;
  assign {FA_cout_2302,FA_out_2302}=FA_out_1424+FA_cout_1485+FA_out_1486;
  assign {FA_cout_2303,FA_out_2303}=FA_out_1425+FA_cout_1486+FA_out_1487;
  assign {FA_cout_2304,FA_out_2304}=FA_out_1426+FA_cout_1487+FA_out_1488;
  assign {FA_cout_2305,FA_out_2305}=FA_out_1427+FA_cout_1488+FA_out_1489;
  assign {FA_cout_2306,FA_out_2306}=FA_out_1428+FA_cout_1489+FA_out_1490;
  assign {FA_cout_2307,FA_out_2307}=FA_out_1429+FA_cout_1490+FA_out_1491;
  assign {FA_cout_2308,FA_out_2308}=FA_out_1430+FA_cout_1491+FA_out_1492;
  assign {FA_cout_2309,FA_out_2309}=FA_out_1431+FA_cout_1492+FA_out_1493;
  assign {FA_cout_2310,FA_out_2310}=FA_out_1432+FA_cout_1493+FA_out_1494;
  assign {FA_cout_2311,FA_out_2311}=FA_out_1433+FA_cout_1494+FA_out_1495;
  assign {FA_cout_2312,FA_out_2312}=FA_out_1434+FA_cout_1495+FA_out_1496;
  assign {FA_cout_2313,FA_out_2313}=FA_out_1435+FA_cout_1496+FA_out_1497;
  assign {FA_cout_2314,FA_out_2314}=FA_out_1436+FA_cout_1497+FA_out_1498;
  assign {FA_cout_2315,FA_out_2315}=FA_out_1437+FA_cout_1498+FA_out_1499;
  assign {FA_cout_2316,FA_out_2316}=FA_out_1438+FA_cout_1499+FA_out_1500;
  assign {FA_cout_2317,FA_out_2317}=FA_out_1439+FA_cout_1500+FA_out_1501;
  assign {FA_cout_2318,FA_out_2318}=FA_out_1440+FA_cout_1501+FA_out_1502;
  assign {FA_cout_2319,FA_out_2319}=FA_out_1441+FA_cout_1502+FA_out_1503;
  assign {FA_cout_2320,FA_out_2320}=FA_out_1442+FA_cout_1503+FA_out_1504;
  assign {FA_cout_2321,FA_out_2321}=FA_out_1443+FA_cout_1504+FA_out_1505;
  assign {FA_cout_2322,FA_out_2322}=FA_out_1444+FA_cout_1505+FA_out_1506;
  assign {FA_cout_2323,FA_out_2323}=FA_out_1446+FA_cout_1506+FA_out_1509;
  assign {FA_cout_2324,FA_out_2324}=FA_cout_1447+FA_out_1449+FA_cout_1507;
  assign {FA_cout_2325,FA_out_2325}=FA_out_1448+FA_cout_1509+FA_out_1512;
  assign {FA_cout_2326,FA_out_2326}=FA_cout_1449+FA_out_1451+FA_cout_1510;
  assign {FA_cout_2327,FA_out_2327}=FA_out_1450+FA_cout_1512+FA_out_1515;
  assign {FA_cout_2328,FA_out_2328}=FA_cout_1451+FA_out_1453+FA_cout_1513;
  assign {FA_cout_2329,FA_out_2329}=FA_out_1452+FA_cout_1515+FA_out_1566;
  assign {FA_cout_2330,FA_out_2330}=FA_cout_1453+FA_out_1508+FA_cout_1516;
  assign {FA_cout_2331,FA_out_2331}=FA_out_1507+FA_cout_1566+FA_out_1570;
  assign {FA_cout_2332,FA_out_2332}=FA_cout_1508+FA_out_1511+FA_cout_1567;
  assign {FA_cout_2333,FA_out_2333}=FA_out_1510+FA_cout_1570+FA_out_1574;
  assign {FA_cout_2334,FA_out_2334}=FA_cout_1511+FA_out_1514+FA_cout_1571;
  assign {FA_cout_2335,FA_out_2335}=FA_out_1513+FA_cout_1574+FA_out_1578;
  assign {FA_cout_2336,FA_out_2336}=FA_cout_1514+FA_out_1517+FA_cout_1575;
  assign {FA_cout_2337,FA_out_2337}=FA_out_1516+FA_cout_1578+FA_out_1582;
  assign {FA_cout_2338,FA_out_2338}=FA_cout_1517+FA_out_1568+FA_cout_1579;
  assign {FA_cout_2339,FA_out_2339}=FA_cout_1518+FA_out_1519+inp_18[0];
  assign {FA_cout_2340,FA_out_2340}=FA_cout_1519+FA_out_1520+HA_out_6;
  assign {FA_cout_2341,FA_out_2341}=FA_cout_1520+FA_out_1521+HA_out_48;
  assign {FA_cout_2342,FA_out_2342}=FA_cout_1521+FA_out_1522+HA_cout_48;
  assign {FA_cout_2343,FA_out_2343}=FA_cout_1522+FA_out_1523+FA_cout_1585;
  assign {FA_cout_2344,FA_out_2344}=FA_cout_1523+FA_out_1524+FA_cout_1586;
  assign {FA_cout_2345,FA_out_2345}=FA_cout_1524+FA_out_1525+FA_cout_1587;
  assign {FA_cout_2346,FA_out_2346}=FA_cout_1525+FA_out_1526+FA_cout_1588;
  assign {FA_cout_2347,FA_out_2347}=FA_cout_1526+FA_out_1527+FA_cout_1589;
  assign {FA_cout_2348,FA_out_2348}=FA_cout_1527+FA_out_1528+FA_cout_1590;
  assign {FA_cout_2349,FA_out_2349}=FA_cout_1528+FA_out_1529+FA_cout_1591;
  assign {FA_cout_2350,FA_out_2350}=FA_cout_1529+FA_out_1530+FA_cout_1592;
  assign {FA_cout_2351,FA_out_2351}=FA_cout_1530+FA_out_1531+FA_cout_1593;
  assign {FA_cout_2352,FA_out_2352}=FA_cout_1531+FA_out_1532+FA_cout_1594;
  assign {FA_cout_2353,FA_out_2353}=FA_cout_1532+FA_out_1533+FA_cout_1595;
  assign {FA_cout_2354,FA_out_2354}=FA_cout_1533+FA_out_1534+FA_cout_1596;
  assign {FA_cout_2355,FA_out_2355}=FA_cout_1534+FA_out_1535+FA_cout_1597;
  assign {FA_cout_2356,FA_out_2356}=FA_cout_1535+FA_out_1536+FA_cout_1598;
  assign {FA_cout_2357,FA_out_2357}=FA_cout_1536+FA_out_1537+FA_cout_1599;
  assign {FA_cout_2358,FA_out_2358}=FA_cout_1537+FA_out_1538+FA_cout_1600;
  assign {FA_cout_2359,FA_out_2359}=FA_cout_1538+FA_out_1539+FA_cout_1601;
  assign {FA_cout_2360,FA_out_2360}=FA_cout_1539+FA_out_1540+FA_cout_1602;
  assign {FA_cout_2361,FA_out_2361}=FA_cout_1540+FA_out_1541+FA_cout_1603;
  assign {FA_cout_2362,FA_out_2362}=FA_cout_1541+FA_out_1542+FA_cout_1604;
  assign {FA_cout_2363,FA_out_2363}=FA_cout_1542+FA_out_1543+FA_cout_1605;
  assign {FA_cout_2364,FA_out_2364}=FA_cout_1543+FA_out_1544+FA_cout_1606;
  assign {FA_cout_2365,FA_out_2365}=FA_cout_1544+FA_out_1545+FA_cout_1607;
  assign {FA_cout_2366,FA_out_2366}=FA_cout_1545+FA_out_1546+FA_cout_1608;
  assign {FA_cout_2367,FA_out_2367}=FA_cout_1546+FA_out_1547+FA_cout_1609;
  assign {FA_cout_2368,FA_out_2368}=FA_cout_1547+FA_out_1548+FA_cout_1610;
  assign {FA_cout_2369,FA_out_2369}=FA_cout_1548+FA_out_1549+FA_cout_1611;
  assign {FA_cout_2370,FA_out_2370}=FA_cout_1549+FA_out_1550+FA_cout_1612;
  assign {FA_cout_2371,FA_out_2371}=FA_cout_1550+FA_out_1551+FA_cout_1613;
  assign {FA_cout_2372,FA_out_2372}=FA_cout_1551+FA_out_1552+FA_cout_1614;
  assign {FA_cout_2373,FA_out_2373}=FA_cout_1552+FA_out_1553+FA_cout_1615;
  assign {FA_cout_2374,FA_out_2374}=FA_cout_1553+FA_out_1554+FA_cout_1616;
  assign {FA_cout_2375,FA_out_2375}=FA_cout_1554+FA_out_1555+FA_cout_1617;
  assign {FA_cout_2376,FA_out_2376}=FA_cout_1555+FA_out_1556+FA_cout_1618;
  assign {FA_cout_2377,FA_out_2377}=FA_cout_1556+FA_out_1557+FA_cout_1619;
  assign {FA_cout_2378,FA_out_2378}=FA_cout_1557+FA_out_1558+FA_cout_1620;
  assign {FA_cout_2379,FA_out_2379}=FA_cout_1558+FA_out_1559+FA_cout_1621;
  assign {FA_cout_2380,FA_out_2380}=FA_cout_1559+FA_out_1560+FA_cout_1622;
  assign {FA_cout_2381,FA_out_2381}=FA_cout_1560+FA_out_1561+FA_cout_1623;
  assign {FA_cout_2382,FA_out_2382}=FA_cout_1561+FA_out_1562+FA_cout_1624;
  assign {FA_cout_2383,FA_out_2383}=FA_cout_1562+FA_out_1563+FA_cout_1625;
  assign {FA_cout_2384,FA_out_2384}=FA_cout_1563+FA_out_1564+FA_cout_1626;
  assign {FA_cout_2385,FA_out_2385}=FA_cout_1564+FA_out_1565+FA_cout_1627;
  assign {FA_cout_2386,FA_out_2386}=FA_cout_1565+FA_out_1569+FA_cout_1628;
  assign {FA_cout_2387,FA_out_2387}=FA_out_1567+FA_cout_1582+FA_out_1630;
  assign {FA_cout_2388,FA_out_2388}=FA_cout_1568+FA_out_1572+FA_cout_1583;
  assign {FA_cout_2389,FA_out_2389}=FA_cout_1569+FA_out_1573+FA_cout_1633;
  assign {FA_cout_2390,FA_out_2390}=FA_out_1571+FA_cout_1630+FA_out_1635;
  assign {FA_cout_2391,FA_out_2391}=FA_cout_1572+FA_out_1576+FA_cout_1631;
  assign {FA_cout_2392,FA_out_2392}=FA_cout_1573+FA_out_1577+FA_cout_1638;
  assign {FA_cout_2393,FA_out_2393}=FA_out_1575+FA_cout_1635+FA_out_1640;
  assign {FA_cout_2394,FA_out_2394}=FA_cout_1576+FA_out_1580+FA_cout_1636;
  assign {FA_cout_2395,FA_out_2395}=FA_cout_1577+FA_out_1581+FA_cout_1643;
  assign {FA_cout_2396,FA_out_2396}=FA_out_1579+FA_cout_1640+FA_out_1645;
  assign {FA_cout_2397,FA_out_2397}=FA_cout_1580+FA_out_1584+FA_cout_1641;
  assign {FA_cout_2398,FA_out_2398}=FA_cout_1581+FA_out_1629+FA_cout_1687;
  assign {FA_cout_2399,FA_out_2399}=FA_out_1583+FA_cout_1645+FA_out_1689;
  assign {FA_cout_2400,FA_out_2400}=FA_cout_1584+FA_out_1632+FA_cout_1646;
  assign {FA_cout_2401,FA_out_2401}=FA_cout_1629+FA_out_1634+FA_cout_1693;
  assign {FA_cout_2402,FA_out_2402}=FA_out_1631+FA_cout_1689+FA_out_1695;
  assign {FA_cout_2403,FA_out_2403}=FA_cout_1632+FA_out_1637+FA_cout_1690;
  assign {FA_cout_2404,FA_out_2404}=FA_out_1589+HA_cout_49+HA_out_50;
  assign {FA_cout_2405,FA_out_2405}=FA_out_1590+HA_cout_50+FA_out_1648;
  assign {FA_cout_2406,FA_out_2406}=FA_out_1591+FA_cout_1648+FA_out_1649;
  assign {FA_cout_2407,FA_out_2407}=FA_out_1592+FA_cout_1649+FA_out_1650;
  assign {FA_cout_2408,FA_out_2408}=FA_out_1593+FA_cout_1650+FA_out_1651;
  assign {FA_cout_2409,FA_out_2409}=FA_out_1594+FA_cout_1651+FA_out_1652;
  assign {FA_cout_2410,FA_out_2410}=FA_out_1595+FA_cout_1652+FA_out_1653;
  assign {FA_cout_2411,FA_out_2411}=FA_out_1596+FA_cout_1653+FA_out_1654;
  assign {FA_cout_2412,FA_out_2412}=FA_out_1597+FA_cout_1654+FA_out_1655;
  assign {FA_cout_2413,FA_out_2413}=FA_out_1598+FA_cout_1655+FA_out_1656;
  assign {FA_cout_2414,FA_out_2414}=FA_out_1599+FA_cout_1656+FA_out_1657;
  assign {FA_cout_2415,FA_out_2415}=FA_out_1600+FA_cout_1657+FA_out_1658;
  assign {FA_cout_2416,FA_out_2416}=FA_out_1601+FA_cout_1658+FA_out_1659;
  assign {FA_cout_2417,FA_out_2417}=FA_out_1602+FA_cout_1659+FA_out_1660;
  assign {FA_cout_2418,FA_out_2418}=FA_out_1603+FA_cout_1660+FA_out_1661;
  assign {FA_cout_2419,FA_out_2419}=FA_out_1604+FA_cout_1661+FA_out_1662;
  assign {FA_cout_2420,FA_out_2420}=FA_out_1605+FA_cout_1662+FA_out_1663;
  assign {FA_cout_2421,FA_out_2421}=FA_out_1606+FA_cout_1663+FA_out_1664;
  assign {FA_cout_2422,FA_out_2422}=FA_out_1607+FA_cout_1664+FA_out_1665;
  assign {FA_cout_2423,FA_out_2423}=FA_out_1608+FA_cout_1665+FA_out_1666;
  assign {FA_cout_2424,FA_out_2424}=FA_out_1609+FA_cout_1666+FA_out_1667;
  assign {FA_cout_2425,FA_out_2425}=FA_out_1610+FA_cout_1667+FA_out_1668;
  assign {FA_cout_2426,FA_out_2426}=FA_out_1611+FA_cout_1668+FA_out_1669;
  assign {FA_cout_2427,FA_out_2427}=FA_out_1612+FA_cout_1669+FA_out_1670;
  assign {FA_cout_2428,FA_out_2428}=FA_out_1613+FA_cout_1670+FA_out_1671;
  assign {FA_cout_2429,FA_out_2429}=FA_out_1614+FA_cout_1671+FA_out_1672;
  assign {FA_cout_2430,FA_out_2430}=FA_out_1615+FA_cout_1672+FA_out_1673;
  assign {FA_cout_2431,FA_out_2431}=FA_out_1616+FA_cout_1673+FA_out_1674;
  assign {FA_cout_2432,FA_out_2432}=FA_out_1617+FA_cout_1674+FA_out_1675;
  assign {FA_cout_2433,FA_out_2433}=FA_out_1618+FA_cout_1675+FA_out_1676;
  assign {FA_cout_2434,FA_out_2434}=FA_out_1619+FA_cout_1676+FA_out_1677;
  assign {FA_cout_2435,FA_out_2435}=FA_out_1620+FA_cout_1677+FA_out_1678;
  assign {FA_cout_2436,FA_out_2436}=FA_out_1621+FA_cout_1678+FA_out_1679;
  assign {FA_cout_2437,FA_out_2437}=FA_out_1622+FA_cout_1679+FA_out_1680;
  assign {FA_cout_2438,FA_out_2438}=FA_out_1623+FA_cout_1680+FA_out_1681;
  assign {FA_cout_2439,FA_out_2439}=FA_out_1624+FA_cout_1681+FA_out_1682;
  assign {FA_cout_2440,FA_out_2440}=FA_out_1625+FA_cout_1682+FA_out_1683;
  assign {FA_cout_2441,FA_out_2441}=FA_out_1626+FA_cout_1683+FA_out_1684;
  assign {FA_cout_2442,FA_out_2442}=FA_out_1627+FA_cout_1684+FA_out_1685;
  assign {FA_cout_2443,FA_out_2443}=FA_out_1628+FA_cout_1685+FA_out_1686;
  assign {FA_cout_2444,FA_out_2444}=FA_out_1633+FA_cout_1686+FA_out_1692;
  assign {FA_cout_2445,FA_out_2445}=FA_cout_1634+FA_out_1639+FA_cout_1699;
  assign {FA_cout_2446,FA_out_2446}=FA_out_1636+FA_cout_1695+FA_out_1701;
  assign {FA_cout_2447,FA_out_2447}=FA_cout_1637+FA_out_1642+FA_cout_1696;
  assign {FA_cout_2448,FA_out_2448}=FA_out_1638+FA_cout_1692+FA_out_1698;
  assign {FA_cout_2449,FA_out_2449}=FA_cout_1639+FA_out_1644+FA_cout_1705;
  assign {FA_cout_2450,FA_out_2450}=FA_out_1641+FA_cout_1701+FA_out_1707;
  assign {FA_cout_2451,FA_out_2451}=FA_cout_1642+FA_out_1647+FA_cout_1702;
  assign {FA_cout_2452,FA_out_2452}=FA_out_1643+FA_cout_1698+FA_out_1704;
  assign {FA_cout_2453,FA_out_2453}=FA_cout_1644+FA_out_1688+FA_cout_1711;
  assign {FA_cout_2454,FA_out_2454}=FA_out_1646+FA_cout_1707+FA_out_1713;
  assign {FA_cout_2455,FA_out_2455}=FA_cout_1647+FA_out_1691+FA_cout_1708;
  assign {FA_cout_2456,FA_out_2456}=FA_out_1687+FA_cout_1704+FA_out_1710;
  assign {FA_cout_2457,FA_out_2457}=FA_cout_1688+FA_out_1694+FA_cout_1752;
  assign {FA_cout_2458,FA_out_2458}=FA_out_1690+FA_cout_1713+FA_out_1754;
  assign {FA_cout_2459,FA_out_2459}=FA_cout_1691+FA_out_1697+FA_cout_1714;
  assign {FA_cout_2460,FA_out_2460}=FA_out_1693+FA_cout_1710+FA_out_1751;
  assign {FA_cout_2461,FA_out_2461}=FA_cout_1694+FA_out_1700+FA_cout_1759;
  assign {FA_cout_2462,FA_out_2462}=FA_out_1696+FA_cout_1754+FA_out_1761;
  assign {FA_cout_2463,FA_out_2463}=FA_cout_1697+FA_out_1703+FA_cout_1755;
  assign {FA_cout_2464,FA_out_2464}=FA_out_1699+FA_cout_1751+FA_out_1758;
  assign {FA_cout_2465,FA_out_2465}=FA_cout_1700+FA_out_1706+FA_cout_1766;
  assign {FA_cout_2466,FA_out_2466}=FA_out_1702+FA_cout_1761+FA_out_1768;
  assign {FA_cout_2467,FA_out_2467}=FA_cout_1703+FA_out_1709+FA_cout_1762;
  assign {FA_cout_2468,FA_out_2468}=FA_out_1705+FA_cout_1758+FA_out_1765;
  assign {FA_cout_2469,FA_out_2469}=FA_cout_1706+FA_out_1712+FA_cout_1773;
  assign {FA_cout_2470,FA_out_2470}=FA_out_1708+FA_cout_1768+FA_out_1775;
  assign {FA_cout_2471,FA_out_2471}=FA_cout_1709+FA_out_1715+FA_cout_1769;
  assign {FA_cout_2472,FA_out_2472}=FA_out_1711+FA_cout_1765+FA_out_1772;
  assign {FA_cout_2473,FA_out_2473}=FA_cout_1712+FA_out_1753+FA_cout_1810;
  assign {FA_cout_2474,FA_out_2474}=FA_out_1714+FA_cout_1775+FA_out_1812;
  assign {FA_cout_2475,FA_out_2475}=FA_cout_1715+FA_out_1756+FA_cout_1776;
  assign {FA_cout_2476,FA_out_2476}=FA_cout_1717+FA_out_1718+FA_out_640;
  assign {FA_cout_2477,FA_out_2477}=FA_cout_1718+FA_out_1719+HA_out_52;
  assign {FA_cout_2478,FA_out_2478}=FA_cout_1719+FA_out_1720+HA_cout_52;
  assign {FA_cout_2479,FA_out_2479}=FA_cout_1720+FA_out_1721+HA_cout_53;
  assign {FA_cout_2480,FA_out_2480}=FA_cout_1721+FA_out_1722+FA_cout_1778;
  assign {FA_cout_2481,FA_out_2481}=FA_cout_1722+FA_out_1723+FA_cout_1779;
  assign {FA_cout_2482,FA_out_2482}=FA_cout_1723+FA_out_1724+FA_cout_1780;
  assign {FA_cout_2483,FA_out_2483}=FA_cout_1724+FA_out_1725+FA_cout_1781;
  assign {FA_cout_2484,FA_out_2484}=FA_cout_1725+FA_out_1726+FA_cout_1782;
  assign {FA_cout_2485,FA_out_2485}=FA_cout_1726+FA_out_1727+FA_cout_1783;
  assign {FA_cout_2486,FA_out_2486}=FA_cout_1727+FA_out_1728+FA_cout_1784;
  assign {FA_cout_2487,FA_out_2487}=FA_cout_1728+FA_out_1729+FA_cout_1785;
  assign {FA_cout_2488,FA_out_2488}=FA_cout_1729+FA_out_1730+FA_cout_1786;
  assign {FA_cout_2489,FA_out_2489}=FA_cout_1730+FA_out_1731+FA_cout_1787;
  assign {FA_cout_2490,FA_out_2490}=FA_cout_1731+FA_out_1732+FA_cout_1788;
  assign {FA_cout_2491,FA_out_2491}=FA_cout_1732+FA_out_1733+FA_cout_1789;
  assign {FA_cout_2492,FA_out_2492}=FA_cout_1733+FA_out_1734+FA_cout_1790;
  assign {FA_cout_2493,FA_out_2493}=FA_cout_1734+FA_out_1735+FA_cout_1791;
  assign {FA_cout_2494,FA_out_2494}=FA_cout_1735+FA_out_1736+FA_cout_1792;
  assign {FA_cout_2495,FA_out_2495}=FA_cout_1736+FA_out_1737+FA_cout_1793;
  assign {FA_cout_2496,FA_out_2496}=FA_cout_1737+FA_out_1738+FA_cout_1794;
  assign {FA_cout_2497,FA_out_2497}=FA_cout_1738+FA_out_1739+FA_cout_1795;
  assign {FA_cout_2498,FA_out_2498}=FA_cout_1739+FA_out_1740+FA_cout_1796;
  assign {FA_cout_2499,FA_out_2499}=FA_cout_1740+FA_out_1741+FA_cout_1797;
  assign {FA_cout_2500,FA_out_2500}=FA_cout_1741+FA_out_1742+FA_cout_1798;
  assign {FA_cout_2501,FA_out_2501}=FA_cout_1742+FA_out_1743+FA_cout_1799;
  assign {FA_cout_2502,FA_out_2502}=FA_cout_1743+FA_out_1744+FA_cout_1800;
  assign {FA_cout_2503,FA_out_2503}=FA_cout_1744+FA_out_1745+FA_cout_1801;
  assign {FA_cout_2504,FA_out_2504}=FA_cout_1745+FA_out_1746+FA_cout_1802;
  assign {FA_cout_2505,FA_out_2505}=FA_cout_1746+FA_out_1747+FA_cout_1803;
  assign {FA_cout_2506,FA_out_2506}=FA_cout_1747+FA_out_1748+FA_cout_1804;
  assign {FA_cout_2507,FA_out_2507}=FA_cout_1748+FA_out_1749+FA_cout_1805;
  assign {FA_cout_2508,FA_out_2508}=FA_cout_1749+FA_out_1750+FA_cout_1806;
  assign {FA_cout_2509,FA_out_2509}=FA_cout_1750+FA_out_1757+FA_cout_1807;
  assign {FA_cout_2510,FA_out_2510}=FA_out_1752+FA_cout_1772+FA_out_1809;
  assign {FA_cout_2511,FA_out_2511}=FA_cout_1753+FA_out_1760+FA_cout_1818;
  assign {FA_cout_2512,FA_out_2512}=FA_out_1755+FA_cout_1812+FA_out_1820;
  assign {FA_cout_2513,FA_out_2513}=FA_cout_1756+FA_out_1763+FA_cout_1813;
  assign {FA_cout_2514,FA_out_2514}=FA_cout_1757+FA_out_1764+FA_cout_1815;
  assign {FA_cout_2515,FA_out_2515}=FA_out_1759+FA_cout_1809+FA_out_1817;
  assign {FA_cout_2516,FA_out_2516}=FA_cout_1760+FA_out_1767+FA_cout_1826;
  assign {FA_cout_2517,FA_out_2517}=FA_out_1762+FA_cout_1820+FA_out_1828;
  assign {FA_cout_2518,FA_out_2518}=FA_cout_1763+FA_out_1770+FA_cout_1821;
  assign {FA_cout_2519,FA_out_2519}=FA_cout_1764+FA_out_1771+FA_cout_1823;
  assign {FA_cout_2520,FA_out_2520}=FA_out_1766+FA_cout_1817+FA_out_1825;
  assign {FA_cout_2521,FA_out_2521}=FA_cout_1767+FA_out_1774+FA_cout_1834;
  assign {FA_cout_2522,FA_out_2522}=FA_out_1769+FA_cout_1828+FA_out_1836;
  assign {FA_cout_2523,FA_out_2523}=FA_cout_1770+FA_out_1777+FA_cout_1829;
  assign {FA_cout_2524,FA_out_2524}=FA_cout_1771+FA_out_1808+FA_cout_1831;
  assign {FA_cout_2525,FA_out_2525}=FA_out_1773+FA_cout_1825+FA_out_1833;
  assign {FA_cout_2526,FA_out_2526}=FA_cout_1774+FA_out_1811+FA_cout_1842;
  assign {FA_cout_2527,FA_out_2527}=FA_out_1776+FA_cout_1836+FA_out_1844;
  assign {FA_cout_2528,FA_out_2528}=FA_cout_1777+FA_out_1814+FA_cout_1837;
  assign {FA_cout_2529,FA_out_2529}=FA_cout_1808+FA_out_1816+FA_cout_1839;
  assign {FA_cout_2530,FA_out_2530}=FA_out_1810+FA_cout_1833+FA_out_1841;
  assign {FA_cout_2531,FA_out_2531}=FA_cout_1811+FA_out_1819+FA_cout_1876;
  assign {FA_cout_2532,FA_out_2532}=FA_out_1813+FA_cout_1844+FA_out_1878;
  assign {FA_cout_2533,FA_out_2533}=FA_cout_1814+FA_out_1822+FA_cout_1845;
  assign {FA_cout_2534,FA_out_2534}=FA_out_1782+HA_cout_54+FA_out_1847;
  assign {FA_cout_2535,FA_out_2535}=FA_out_1783+FA_cout_1847+FA_out_1848;
  assign {FA_cout_2536,FA_out_2536}=FA_out_1784+FA_cout_1848+FA_out_1849;
  assign {FA_cout_2537,FA_out_2537}=FA_out_1785+FA_cout_1849+FA_out_1850;
  assign {FA_cout_2538,FA_out_2538}=FA_out_1786+FA_cout_1850+FA_out_1851;
  assign {FA_cout_2539,FA_out_2539}=FA_out_1787+FA_cout_1851+FA_out_1852;
  assign {FA_cout_2540,FA_out_2540}=FA_out_1788+FA_cout_1852+FA_out_1853;
  assign {FA_cout_2541,FA_out_2541}=FA_out_1789+FA_cout_1853+FA_out_1854;
  assign {FA_cout_2542,FA_out_2542}=FA_out_1790+FA_cout_1854+FA_out_1855;
  assign {FA_cout_2543,FA_out_2543}=FA_out_1791+FA_cout_1855+FA_out_1856;
  assign {FA_cout_2544,FA_out_2544}=FA_out_1792+FA_cout_1856+FA_out_1857;
  assign {FA_cout_2545,FA_out_2545}=FA_out_1793+FA_cout_1857+FA_out_1858;
  assign {FA_cout_2546,FA_out_2546}=FA_out_1794+FA_cout_1858+FA_out_1859;
  assign {FA_cout_2547,FA_out_2547}=FA_out_1795+FA_cout_1859+FA_out_1860;
  assign {FA_cout_2548,FA_out_2548}=FA_out_1796+FA_cout_1860+FA_out_1861;
  assign {FA_cout_2549,FA_out_2549}=FA_out_1797+FA_cout_1861+FA_out_1862;
  assign {FA_cout_2550,FA_out_2550}=FA_out_1798+FA_cout_1862+FA_out_1863;
  assign {FA_cout_2551,FA_out_2551}=FA_out_1799+FA_cout_1863+FA_out_1864;
  assign {FA_cout_2552,FA_out_2552}=FA_out_1800+FA_cout_1864+FA_out_1865;
  assign {FA_cout_2553,FA_out_2553}=FA_out_1801+FA_cout_1865+FA_out_1866;
  assign {FA_cout_2554,FA_out_2554}=FA_out_1802+FA_cout_1866+FA_out_1867;
  assign {FA_cout_2555,FA_out_2555}=FA_out_1803+FA_cout_1867+FA_out_1868;
  assign {FA_cout_2556,FA_out_2556}=FA_out_1804+FA_cout_1868+FA_out_1869;
  assign {FA_cout_2557,FA_out_2557}=FA_out_1805+FA_cout_1869+FA_out_1870;
  assign {FA_cout_2558,FA_out_2558}=FA_out_1806+FA_cout_1870+FA_out_1871;
  assign {FA_cout_2559,FA_out_2559}=FA_out_1807+FA_cout_1871+FA_out_1872;
  assign {FA_cout_2560,FA_out_2560}=FA_out_1815+FA_cout_1872+FA_out_1881;
  assign {FA_cout_2561,FA_out_2561}=FA_cout_1816+FA_out_1824+FA_cout_1873;
  assign {FA_cout_2562,FA_out_2562}=FA_out_1818+FA_cout_1841+FA_out_1875;
  assign {FA_cout_2563,FA_out_2563}=FA_cout_1819+FA_out_1827+FA_cout_1885;
  assign {FA_cout_2564,FA_out_2564}=FA_out_1821+FA_cout_1878+FA_out_1887;
  assign {FA_cout_2565,FA_out_2565}=FA_cout_1822+FA_out_1830+FA_cout_1879;
  assign {FA_cout_2566,FA_out_2566}=FA_out_1823+FA_cout_1881+FA_out_1890;
  assign {FA_cout_2567,FA_out_2567}=FA_cout_1824+FA_out_1832+FA_cout_1882;
  assign {FA_cout_2568,FA_out_2568}=FA_out_1826+FA_cout_1875+FA_out_1884;
  assign {FA_cout_2569,FA_out_2569}=FA_cout_1827+FA_out_1835+FA_cout_1894;
  assign {FA_cout_2570,FA_out_2570}=FA_out_1829+FA_cout_1887+FA_out_1896;
  assign {FA_cout_2571,FA_out_2571}=FA_cout_1830+FA_out_1838+FA_cout_1888;
  assign {FA_cout_2572,FA_out_2572}=FA_out_1831+FA_cout_1890+FA_out_1899;
  assign {FA_cout_2573,FA_out_2573}=FA_cout_1832+FA_out_1840+FA_cout_1891;
  assign {FA_cout_2574,FA_out_2574}=FA_out_1834+FA_cout_1884+FA_out_1893;
  assign {FA_cout_2575,FA_out_2575}=FA_cout_1835+FA_out_1843+FA_cout_1903;
  assign {FA_cout_2576,FA_out_2576}=FA_out_1837+FA_cout_1896+FA_out_1905;
  assign {FA_cout_2577,FA_out_2577}=FA_cout_1838+FA_out_1846+FA_cout_1897;
  assign {FA_cout_2578,FA_out_2578}=FA_out_1839+FA_cout_1899+FA_out_1929;
  assign {FA_cout_2579,FA_out_2579}=FA_cout_1840+FA_out_1874+FA_cout_1900;
  assign {FA_cout_2580,FA_out_2580}=FA_out_1842+FA_cout_1893+FA_out_1902;
  assign {FA_cout_2581,FA_out_2581}=FA_cout_1843+FA_out_1877+FA_cout_1933;
  assign {FA_cout_2582,FA_out_2582}=FA_out_1845+FA_cout_1905+FA_out_1935;
  assign {FA_cout_2583,FA_out_2583}=FA_cout_1846+FA_out_1880+FA_cout_1906;
  assign {FA_cout_2584,FA_out_2584}=FA_out_1873+FA_cout_1929+FA_out_1939;
  assign {FA_cout_2585,FA_out_2585}=FA_cout_1874+FA_out_1883+FA_cout_1930;
  assign {FA_cout_2586,FA_out_2586}=FA_out_1876+FA_cout_1902+FA_out_1932;
  assign {FA_cout_2587,FA_out_2587}=FA_cout_1877+FA_out_1886+FA_cout_1943;
  assign {FA_cout_2588,FA_out_2588}=FA_out_1879+FA_cout_1935+FA_out_1945;
  assign {FA_cout_2589,FA_out_2589}=FA_cout_1880+FA_out_1889+FA_cout_1936;
  assign {FA_cout_2590,FA_out_2590}=FA_out_1882+FA_cout_1939+FA_out_1949;
  assign {FA_cout_2591,FA_out_2591}=FA_cout_1883+FA_out_1892+FA_cout_1940;
  assign {FA_cout_2592,FA_out_2592}=FA_out_1885+FA_cout_1932+FA_out_1942;
  assign {FA_cout_2593,FA_out_2593}=FA_cout_1886+FA_out_1895+FA_cout_1953;
  assign {FA_cout_2594,FA_out_2594}=FA_out_1888+FA_cout_1945+FA_out_1955;
  assign {FA_cout_2595,FA_out_2595}=FA_cout_1889+FA_out_1898+FA_cout_1946;
  assign {FA_cout_2596,FA_out_2596}=FA_out_1891+FA_cout_1949+FA_out_1959;
  assign {FA_cout_2597,FA_out_2597}=FA_cout_1892+FA_out_1901+FA_cout_1950;
  assign {FA_cout_2598,FA_out_2598}=FA_out_1894+FA_cout_1942+FA_out_1952;
  assign {FA_cout_2599,FA_out_2599}=FA_cout_1895+FA_out_1904+FA_cout_1963;
  assign {FA_cout_2600,FA_out_2600}=FA_out_1897+FA_cout_1955+FA_out_1965;
  assign {FA_cout_2601,FA_out_2601}=FA_cout_1898+FA_out_1907+FA_cout_1956;
  assign {FA_cout_2602,FA_out_2602}=FA_out_1900+FA_cout_1959+FA_out_1969;
  assign {FA_cout_2603,FA_out_2603}=FA_cout_1901+FA_out_1931+FA_cout_1960;
  assign {FA_cout_2604,FA_out_2604}=FA_out_1903+FA_cout_1952+FA_out_1962;
  assign {FA_cout_2605,FA_out_2605}=FA_cout_1904+FA_out_1934+FA_cout_1973;
  assign {FA_cout_2606,FA_out_2606}=FA_out_1906+FA_cout_1965+FA_out_1975;
  assign {FA_cout_2607,FA_out_2607}=FA_cout_1907+FA_out_1937+FA_cout_1966;
  assign {FA_cout_2608,FA_out_2608}=FA_cout_1908+FA_out_1909+inp_45[0];
  assign {FA_cout_2609,FA_out_2609}=FA_cout_1909+FA_out_1910+HA_out_15;
  assign {FA_cout_2610,FA_out_2610}=FA_cout_1910+FA_out_1911+HA_out_57;
  assign {FA_cout_2611,FA_out_2611}=FA_cout_1911+FA_out_1912+HA_cout_57;
  assign {FA_cout_2612,FA_out_2612}=FA_cout_1912+FA_out_1913+FA_cout_1978;
  assign {FA_cout_2613,FA_out_2613}=FA_cout_1913+FA_out_1914+FA_cout_1979;
  assign {FA_cout_2614,FA_out_2614}=FA_cout_1914+FA_out_1915+FA_cout_1980;
  assign {FA_cout_2615,FA_out_2615}=FA_cout_1915+FA_out_1916+FA_cout_1981;
  assign {FA_cout_2616,FA_out_2616}=FA_cout_1916+FA_out_1917+FA_cout_1982;
  assign {FA_cout_2617,FA_out_2617}=FA_cout_1917+FA_out_1918+FA_cout_1983;
  assign {FA_cout_2618,FA_out_2618}=FA_cout_1918+FA_out_1919+FA_cout_1984;
  assign {FA_cout_2619,FA_out_2619}=FA_cout_1919+FA_out_1920+FA_cout_1985;
  assign {FA_cout_2620,FA_out_2620}=FA_cout_1920+FA_out_1921+FA_cout_1986;
  assign {FA_cout_2621,FA_out_2621}=FA_cout_1921+FA_out_1922+FA_cout_1987;
  assign {FA_cout_2622,FA_out_2622}=FA_cout_1922+FA_out_1923+FA_cout_1988;
  assign {FA_cout_2623,FA_out_2623}=FA_cout_1923+FA_out_1924+FA_cout_1989;
  assign {FA_cout_2624,FA_out_2624}=FA_cout_1924+FA_out_1925+FA_cout_1990;
  assign {FA_cout_2625,FA_out_2625}=FA_cout_1925+FA_out_1926+FA_cout_1991;
  assign {FA_cout_2626,FA_out_2626}=FA_cout_1926+FA_out_1927+FA_cout_1992;
  assign {FA_cout_2627,FA_out_2627}=FA_cout_1927+FA_out_1928+FA_cout_1993;
  assign {FA_cout_2628,FA_out_2628}=FA_cout_1928+FA_out_1938+FA_cout_1994;
  assign {FA_cout_2629,FA_out_2629}=FA_out_1930+FA_cout_1969+FA_out_1996;
  assign {FA_cout_2630,FA_out_2630}=FA_cout_1931+FA_out_1941+FA_cout_1970;
  assign {FA_cout_2631,FA_out_2631}=FA_out_1933+FA_cout_1962+FA_out_1972;
  assign {FA_cout_2632,FA_out_2632}=FA_cout_1934+FA_out_1944+FA_cout_2000;
  assign {FA_cout_2633,FA_out_2633}=FA_out_1936+FA_cout_1975+FA_out_2002;
  assign {FA_cout_2634,FA_out_2634}=FA_cout_1937+FA_out_1947+FA_cout_1976;
  assign {FA_cout_2635,FA_out_2635}=FA_cout_1938+FA_out_1948+FA_cout_2005;
  assign {FA_cout_2636,FA_out_2636}=FA_out_1940+FA_cout_1996+FA_out_2007;
  assign {FA_cout_2637,FA_out_2637}=FA_cout_1941+FA_out_1951+FA_cout_1997;
  assign {FA_cout_2638,FA_out_2638}=FA_out_1943+FA_cout_1972+FA_out_1999;
  assign {FA_cout_2639,FA_out_2639}=FA_cout_1944+FA_out_1954+FA_cout_2011;
  assign {FA_cout_2640,FA_out_2640}=FA_out_1946+FA_cout_2002+FA_out_2013;
  assign {FA_cout_2641,FA_out_2641}=FA_cout_1947+FA_out_1957+FA_cout_2003;
  assign {FA_cout_2642,FA_out_2642}=FA_cout_1948+FA_out_1958+FA_cout_2016;
  assign {FA_cout_2643,FA_out_2643}=FA_out_1950+FA_cout_2007+FA_out_2018;
  assign {FA_cout_2644,FA_out_2644}=FA_cout_1951+FA_out_1961+FA_cout_2008;
  assign {FA_cout_2645,FA_out_2645}=FA_out_1953+FA_cout_1999+FA_out_2010;
  assign {FA_cout_2646,FA_out_2646}=FA_cout_1954+FA_out_1964+FA_cout_2022;
  assign {FA_cout_2647,FA_out_2647}=FA_out_1956+FA_cout_2013+FA_out_2024;
  assign {FA_cout_2648,FA_out_2648}=FA_cout_1957+FA_out_1967+FA_cout_2014;
  assign {FA_cout_2649,FA_out_2649}=FA_cout_1958+FA_out_1968+FA_cout_2027;
  assign {FA_cout_2650,FA_out_2650}=FA_out_1960+FA_cout_2018+FA_out_2029;
  assign {FA_cout_2651,FA_out_2651}=FA_cout_1961+FA_out_1971+FA_cout_2019;
  assign {FA_cout_2652,FA_out_2652}=FA_out_1963+FA_cout_2010+FA_out_2021;
  assign {FA_cout_2653,FA_out_2653}=FA_cout_1964+FA_out_1974+FA_cout_2033;
  assign {FA_cout_2654,FA_out_2654}=FA_out_1966+FA_cout_2024+FA_out_2035;
  assign {FA_cout_2655,FA_out_2655}=FA_cout_1967+FA_out_1977+FA_cout_2025;
  assign {FA_cout_2656,FA_out_2656}=FA_cout_1968+FA_out_1995+FA_cout_2050;
  assign {FA_cout_2657,FA_out_2657}=FA_out_1970+FA_cout_2029+FA_out_2052;
  assign {FA_cout_2658,FA_out_2658}=FA_cout_1971+FA_out_1998+FA_cout_2030;
  assign {FA_cout_2659,FA_out_2659}=FA_out_1973+FA_cout_2021+FA_out_2032;
  assign {FA_cout_2660,FA_out_2660}=FA_cout_1974+FA_out_2001+FA_cout_2056;
  assign {FA_cout_2661,FA_out_2661}=FA_out_1976+FA_cout_2035+FA_out_2058;
  assign {FA_cout_2662,FA_out_2662}=FA_cout_1977+FA_out_2004+FA_cout_2036;
  assign {FA_cout_2663,FA_out_2663}=FA_cout_1995+FA_out_2006+FA_cout_2062;
  assign {FA_cout_2664,FA_out_2664}=FA_out_1997+FA_cout_2052+FA_out_2064;
  assign {FA_cout_2665,FA_out_2665}=FA_cout_1998+FA_out_2009+FA_cout_2053;
  assign {FA_cout_2666,FA_out_2666}=FA_out_2000+FA_cout_2032+FA_out_2055;
  assign {FA_cout_2667,FA_out_2667}=FA_cout_2001+FA_out_2012+FA_cout_2068;
  assign {FA_cout_2668,FA_out_2668}=FA_out_2003+FA_cout_2058+FA_out_2070;
  assign {FA_cout_2669,FA_out_2669}=FA_cout_2004+FA_out_2015+FA_cout_2059;
  assign {FA_cout_2670,FA_out_2670}=FA_out_1982+HA_cout_58+HA_out_59;
  assign {FA_cout_2671,FA_out_2671}=FA_out_1983+HA_cout_59+FA_out_2038;
  assign {FA_cout_2672,FA_out_2672}=FA_out_1984+FA_cout_2038+FA_out_2039;
  assign {FA_cout_2673,FA_out_2673}=FA_out_1985+FA_cout_2039+FA_out_2040;
  assign {FA_cout_2674,FA_out_2674}=FA_out_1986+FA_cout_2040+FA_out_2041;
  assign {FA_cout_2675,FA_out_2675}=FA_out_1987+FA_cout_2041+FA_out_2042;
  assign {FA_cout_2676,FA_out_2676}=FA_out_1988+FA_cout_2042+FA_out_2043;
  assign {FA_cout_2677,FA_out_2677}=FA_out_1989+FA_cout_2043+FA_out_2044;
  assign {FA_cout_2678,FA_out_2678}=FA_out_1990+FA_cout_2044+FA_out_2045;
  assign {FA_cout_2679,FA_out_2679}=FA_out_1991+FA_cout_2045+FA_out_2046;
  assign {FA_cout_2680,FA_out_2680}=FA_out_1992+FA_cout_2046+FA_out_2047;
  assign {FA_cout_2681,FA_out_2681}=FA_out_1993+FA_cout_2047+FA_out_2048;
  assign {FA_cout_2682,FA_out_2682}=FA_out_1994+FA_cout_2048+FA_out_2049;
  assign {FA_cout_2683,FA_out_2683}=FA_out_2005+FA_cout_2049+FA_out_2061;
  assign {FA_cout_2684,FA_out_2684}=FA_cout_2006+FA_out_2017+FA_cout_2074;
  assign {FA_cout_2685,FA_out_2685}=FA_out_2008+FA_cout_2064+FA_out_2076;
  assign {FA_cout_2686,FA_out_2686}=FA_cout_2009+FA_out_2020+FA_cout_2065;
  assign {FA_cout_2687,FA_out_2687}=FA_out_2011+FA_cout_2055+FA_out_2067;
  assign {FA_cout_2688,FA_out_2688}=FA_cout_2012+FA_out_2023+FA_cout_2080;
  assign {FA_cout_2689,FA_out_2689}=FA_out_2014+FA_cout_2070+FA_out_2082;
  assign {FA_cout_2690,FA_out_2690}=FA_cout_2015+FA_out_2026+FA_cout_2071;
  assign {FA_cout_2691,FA_out_2691}=FA_out_2016+FA_cout_2061+FA_out_2073;
  assign {FA_cout_2692,FA_out_2692}=FA_cout_2017+FA_out_2028+FA_cout_2086;
  assign {FA_cout_2693,FA_out_2693}=FA_out_2019+FA_cout_2076+FA_out_2088;
  assign {FA_cout_2694,FA_out_2694}=FA_cout_2020+FA_out_2031+FA_cout_2077;
  assign {FA_cout_2695,FA_out_2695}=FA_out_2022+FA_cout_2067+FA_out_2079;
  assign {FA_cout_2696,FA_out_2696}=FA_cout_2023+FA_out_2034+FA_cout_2092;
  assign {FA_cout_2697,FA_out_2697}=FA_out_2025+FA_cout_2082+FA_out_2094;
  assign {FA_cout_2698,FA_out_2698}=FA_cout_2026+FA_out_2037+FA_cout_2083;
  assign {FA_cout_2699,FA_out_2699}=FA_out_2027+FA_cout_2073+FA_out_2085;
  assign {FA_cout_2700,FA_out_2700}=FA_cout_2028+FA_out_2051+FA_cout_2098;
  assign {FA_cout_2701,FA_out_2701}=FA_out_2030+FA_cout_2088+FA_out_2100;
  assign {FA_cout_2702,FA_out_2702}=FA_cout_2031+FA_out_2054+FA_cout_2089;
  assign {FA_cout_2703,FA_out_2703}=FA_out_2033+FA_cout_2079+FA_out_2091;
  assign {FA_cout_2704,FA_out_2704}=FA_cout_2034+FA_out_2057+FA_cout_2104;
  assign {FA_cout_2705,FA_out_2705}=FA_out_2036+FA_cout_2094+FA_out_2106;
  assign {FA_cout_2706,FA_out_2706}=FA_cout_2037+FA_out_2060+FA_cout_2095;
  assign {FA_cout_2707,FA_out_2707}=FA_out_2050+FA_cout_2085+FA_out_2097;
  assign {FA_cout_2708,FA_out_2708}=FA_cout_2051+FA_out_2063+FA_cout_2118;
  assign {FA_cout_2709,FA_out_2709}=FA_out_2053+FA_cout_2100+FA_out_2120;
  assign {FA_cout_2710,FA_out_2710}=FA_cout_2054+FA_out_2066+FA_cout_2101;
  assign {FA_cout_2711,FA_out_2711}=FA_out_2056+FA_cout_2091+FA_out_2103;
  assign {FA_cout_2712,FA_out_2712}=FA_cout_2057+FA_out_2069+FA_cout_2124;
  assign {FA_cout_2713,FA_out_2713}=FA_out_2059+FA_cout_2106+FA_out_2126;
  assign {FA_cout_2714,FA_out_2714}=FA_cout_2060+FA_out_2072+FA_cout_2107;
  assign {FA_cout_2715,FA_out_2715}=FA_out_2062+FA_cout_2097+FA_out_2117;
  assign {FA_cout_2716,FA_out_2716}=FA_cout_2063+FA_out_2075+FA_cout_2131;
  assign {FA_cout_2717,FA_out_2717}=FA_out_2065+FA_cout_2120+FA_out_2133;
  assign {FA_cout_2718,FA_out_2718}=FA_cout_2066+FA_out_2078+FA_cout_2121;
  assign {FA_cout_2719,FA_out_2719}=FA_out_2068+FA_cout_2103+FA_out_2123;
  assign {FA_cout_2720,FA_out_2720}=FA_cout_2069+FA_out_2081+FA_cout_2137;
  assign {FA_cout_2721,FA_out_2721}=FA_out_2071+FA_cout_2126+FA_out_2139;
  assign {FA_cout_2722,FA_out_2722}=FA_cout_2072+FA_out_2084+FA_cout_2127;
  assign {FA_cout_2723,FA_out_2723}=FA_out_2074+FA_cout_2117+FA_out_2130;
  assign {FA_cout_2724,FA_out_2724}=FA_cout_2075+FA_out_2087+FA_cout_2144;
  assign {FA_cout_2725,FA_out_2725}=FA_out_2077+FA_cout_2133+FA_out_2146;
  assign {FA_cout_2726,FA_out_2726}=FA_cout_2078+FA_out_2090+FA_cout_2134;
  assign {FA_cout_2727,FA_out_2727}=FA_out_2080+FA_cout_2123+FA_out_2136;
  assign {FA_cout_2728,FA_out_2728}=FA_cout_2081+FA_out_2093+FA_cout_2150;
  assign {FA_cout_2729,FA_out_2729}=FA_out_2083+FA_cout_2139+FA_out_2152;
  assign {FA_cout_2730,FA_out_2730}=FA_cout_2084+FA_out_2096+FA_cout_2140;
  assign {FA_cout_2731,FA_out_2731}=FA_out_2086+FA_cout_2130+FA_out_2143;
  assign {FA_cout_2732,FA_out_2732}=FA_cout_2087+FA_out_2099+FA_cout_2157;
  assign {FA_cout_2733,FA_out_2733}=FA_out_2089+FA_cout_2146+FA_out_2159;
  assign {FA_cout_2734,FA_out_2734}=FA_cout_2090+FA_out_2102+FA_cout_2147;
  assign {FA_cout_2735,FA_out_2735}=FA_out_2092+FA_cout_2136+FA_out_2149;
  assign {FA_cout_2736,FA_out_2736}=FA_cout_2093+FA_out_2105+FA_cout_2163;
  assign {FA_cout_2737,FA_out_2737}=FA_out_2095+FA_cout_2152+FA_out_2165;
  assign {FA_cout_2738,FA_out_2738}=FA_cout_2096+FA_out_2108+FA_cout_2153;
  assign {FA_cout_2739,FA_out_2739}=FA_out_2098+FA_cout_2143+FA_out_2156;
  assign {FA_cout_2740,FA_out_2740}=FA_cout_2099+FA_out_2119+FA_cout_2173;
  assign {FA_cout_2741,FA_out_2741}=FA_out_2101+FA_cout_2159+FA_out_2175;
  assign {FA_cout_2742,FA_out_2742}=FA_cout_2102+FA_out_2122+FA_cout_2160;
  assign {FA_cout_2743,FA_out_2743}=FA_out_2104+FA_cout_2149+FA_out_2162;
  assign {FA_cout_2744,FA_out_2744}=FA_cout_2105+FA_out_2125+FA_cout_2179;
  assign {FA_cout_2745,FA_out_2745}=FA_out_2107+FA_cout_2165+FA_out_2181;
  assign {FA_cout_2746,FA_out_2746}=FA_cout_2108+FA_out_2128+FA_cout_2166;
  assign {FA_cout_2747,FA_out_2747}=FA_cout_2110+FA_out_2111+FA_out_1216;
  assign {FA_cout_2748,FA_out_2748}=FA_cout_2111+FA_out_2112+HA_out_61;
  assign {FA_cout_2749,FA_out_2749}=FA_cout_2112+FA_out_2113+HA_cout_61;
  assign {FA_cout_2750,FA_out_2750}=FA_cout_2113+FA_out_2114+HA_cout_62;
  assign {FA_cout_2751,FA_out_2751}=FA_cout_2114+FA_out_2115+FA_cout_2168;
  assign {FA_cout_2752,FA_out_2752}=FA_cout_2115+FA_out_2116+FA_cout_2169;
  assign {FA_cout_2753,FA_out_2753}=FA_cout_2116+FA_out_2129+FA_cout_2170;
  assign {FA_cout_2754,FA_out_2754}=FA_out_2118+FA_cout_2156+FA_out_2172;
  assign {FA_cout_2755,FA_out_2755}=FA_cout_2119+FA_out_2132+FA_cout_2187;
  assign {FA_cout_2756,FA_out_2756}=FA_out_2121+FA_cout_2175+FA_out_2189;
  assign {FA_cout_2757,FA_out_2757}=FA_cout_2122+FA_out_2135+FA_cout_2176;
  assign {FA_cout_2758,FA_out_2758}=FA_out_2124+FA_cout_2162+FA_out_2178;
  assign {FA_cout_2759,FA_out_2759}=FA_cout_2125+FA_out_2138+FA_cout_2193;
  assign {FA_cout_2760,FA_out_2760}=FA_out_2127+FA_cout_2181+FA_out_2195;
  assign {FA_cout_2761,FA_out_2761}=FA_cout_2128+FA_out_2141+FA_cout_2182;
  assign {FA_cout_2762,FA_out_2762}=FA_cout_2129+FA_out_2142+FA_cout_2184;
  assign {FA_cout_2763,FA_out_2763}=FA_out_2131+FA_cout_2172+FA_out_2186;
  assign {FA_cout_2764,FA_out_2764}=FA_cout_2132+FA_out_2145+HA_cout_64;
  assign {FA_cout_2765,FA_out_2765}=FA_out_2134+FA_cout_2189+HA_out_65;
  assign {FA_cout_2766,FA_out_2766}=FA_cout_2135+FA_out_2148+FA_cout_2190;
  assign {FA_cout_2767,FA_out_2767}=FA_out_2137+FA_cout_2178+FA_out_2192;
  assign {FA_cout_2768,FA_out_2768}=FA_cout_2138+FA_out_2151+HA_cout_67;
  assign {FA_cout_2769,FA_out_2769}=FA_out_2140+FA_cout_2195+HA_out_68;
  assign {FA_cout_2770,FA_out_2770}=FA_cout_2141+FA_out_2154+FA_cout_2196;
  assign {FA_cout_2771,FA_out_2771}=FA_cout_2142+FA_out_2155+FA_cout_2198;
  assign {FA_cout_2772,FA_out_2772}=FA_out_2144+FA_cout_2186+FA_out_2199;
  assign {FA_cout_2773,FA_out_2773}=FA_cout_2145+FA_out_2158+HA_cout_71;
  assign {FA_cout_2774,FA_out_2774}=FA_out_2147+HA_cout_65+HA_out_72;
  assign {FA_cout_2775,FA_out_2775}=FA_cout_2148+FA_out_2161+FA_cout_2201;
  assign {FA_cout_2776,FA_out_2776}=FA_out_2150+FA_cout_2192+FA_out_2202;
  assign {FA_cout_2777,FA_out_2777}=FA_cout_2151+FA_out_2164+HA_cout_74;
  assign {FA_cout_2778,FA_out_2778}=FA_out_2153+HA_cout_68+HA_out_75;
  assign {FA_cout_2779,FA_out_2779}=FA_cout_2154+FA_out_2167+FA_cout_2204;
  assign {FA_cout_2780,FA_out_2780}=FA_cout_2155+FA_out_2171+HA_out_22;
  assign {FA_cout_2781,FA_out_2781}=FA_out_2157+FA_cout_2199+FA_out_1306;
  assign {FA_cout_2782,FA_out_2782}=FA_cout_2158+FA_out_2174+HA_cout_78;
  assign {FA_cout_2783,FA_out_2783}=FA_out_2160+HA_cout_72+HA_out_79;
  assign {FA_cout_2784,FA_out_2784}=FA_cout_2161+FA_out_2177+HA_out_31;
  assign {FA_cout_2785,FA_out_2785}=FA_out_2163+FA_cout_2202+FA_out_1315;
  assign {FA_cout_2786,FA_out_2786}=FA_cout_2164+FA_out_2180+HA_cout_81;
  assign {FA_cout_2787,FA_out_2787}=FA_out_2166+HA_cout_75+HA_out_82;
  assign {FA_cout_2788,FA_out_2788}=FA_cout_2167+FA_out_2183+HA_out_40;
  assign {FA_cout_2789,FA_out_2789}=FA_cout_2171+FA_out_2185+inp_63[6];
  assign {FA_cout_2790,FA_out_2790}=FA_cout_2177+FA_out_2191+inp_63[33];
  assign {FA_cout_2791,FA_out_2791}=FA_cout_2183+FA_out_2197+inp_63[60];
  assign {FA_cout_2792,FA_out_2792}=REGS_7+REGS_70+REGS_137;
  assign {FA_cout_2793,FA_out_2793}=REGS_8+REGS_71+REGS_138;
  assign {FA_cout_2794,FA_out_2794}=REGS_9+REGS_72+REGS_139;
  assign {FA_cout_2795,FA_out_2795}=REGS_10+REGS_73+REGS_140;
  assign {FA_cout_2796,FA_out_2796}=REGS_11+REGS_74+REGS_141;
  assign {FA_cout_2797,FA_out_2797}=REGS_12+REGS_75+REGS_142;
  assign {FA_cout_2798,FA_out_2798}=REGS_13+REGS_76+REGS_143;
  assign {FA_cout_2799,FA_out_2799}=REGS_14+REGS_77+REGS_144;
  assign {FA_cout_2800,FA_out_2800}=REGS_15+REGS_78+REGS_145;
  assign {FA_cout_2801,FA_out_2801}=REGS_16+REGS_79+REGS_146;
  assign {FA_cout_2802,FA_out_2802}=REGS_17+REGS_80+REGS_147;
  assign {FA_cout_2803,FA_out_2803}=REGS_18+REGS_81+REGS_148;
  assign {FA_cout_2804,FA_out_2804}=REGS_19+REGS_82+REGS_149;
  assign {FA_cout_2805,FA_out_2805}=REGS_20+REGS_83+REGS_150;
  assign {FA_cout_2806,FA_out_2806}=REGS_21+REGS_84+REGS_151;
  assign {FA_cout_2807,FA_out_2807}=REGS_22+REGS_85+REGS_152;
  assign {FA_cout_2808,FA_out_2808}=REGS_23+REGS_86+REGS_153;
  assign {FA_cout_2809,FA_out_2809}=REGS_24+REGS_87+REGS_154;
  assign {FA_cout_2810,FA_out_2810}=REGS_25+REGS_88+REGS_155;
  assign {FA_cout_2811,FA_out_2811}=REGS_26+REGS_89+REGS_156;
  assign {FA_cout_2812,FA_out_2812}=REGS_27+REGS_90+REGS_157;
  assign {FA_cout_2813,FA_out_2813}=REGS_28+REGS_91+REGS_158;
  assign {FA_cout_2814,FA_out_2814}=REGS_29+REGS_92+REGS_159;
  assign {FA_cout_2815,FA_out_2815}=REGS_30+REGS_93+REGS_160;
  assign {FA_cout_2816,FA_out_2816}=REGS_31+REGS_94+REGS_161;
  assign {FA_cout_2817,FA_out_2817}=REGS_32+REGS_95+REGS_162;
  assign {FA_cout_2818,FA_out_2818}=REGS_33+REGS_96+REGS_163;
  assign {FA_cout_2819,FA_out_2819}=REGS_34+REGS_97+REGS_164;
  assign {FA_cout_2820,FA_out_2820}=REGS_35+REGS_98+REGS_165;
  assign {FA_cout_2821,FA_out_2821}=REGS_36+REGS_99+REGS_166;
  assign {FA_cout_2822,FA_out_2822}=REGS_37+REGS_100+REGS_167;
  assign {FA_cout_2823,FA_out_2823}=REGS_38+REGS_101+REGS_168;
  assign {FA_cout_2824,FA_out_2824}=REGS_39+REGS_102+REGS_169;
  assign {FA_cout_2825,FA_out_2825}=REGS_40+REGS_103+REGS_170;
  assign {FA_cout_2826,FA_out_2826}=REGS_41+REGS_104+REGS_171;
  assign {FA_cout_2827,FA_out_2827}=REGS_42+REGS_105+REGS_172;
  assign {FA_cout_2828,FA_out_2828}=REGS_43+REGS_106+REGS_173;
  assign {FA_cout_2829,FA_out_2829}=REGS_44+REGS_107+REGS_174;
  assign {FA_cout_2830,FA_out_2830}=REGS_45+REGS_108+REGS_175;
  assign {FA_cout_2831,FA_out_2831}=REGS_46+REGS_109+REGS_176;
  assign {FA_cout_2832,FA_out_2832}=REGS_47+REGS_110+REGS_177;
  assign {FA_cout_2833,FA_out_2833}=REGS_48+REGS_111+REGS_178;
  assign {FA_cout_2834,FA_out_2834}=REGS_49+REGS_112+REGS_179;
  assign {FA_cout_2835,FA_out_2835}=REGS_50+REGS_113+REGS_180;
  assign {FA_cout_2836,FA_out_2836}=REGS_51+REGS_114+REGS_181;
  assign {FA_cout_2837,FA_out_2837}=REGS_52+REGS_115+REGS_182;
  assign {FA_cout_2838,FA_out_2838}=REGS_53+REGS_116+REGS_183;
  assign {FA_cout_2839,FA_out_2839}=REGS_54+REGS_117+REGS_184;
  assign {FA_cout_2840,FA_out_2840}=REGS_55+REGS_118+REGS_185;
  assign {FA_cout_2841,FA_out_2841}=REGS_56+REGS_119+REGS_186;
  assign {FA_cout_2842,FA_out_2842}=REGS_57+REGS_120+REGS_187;
  assign {FA_cout_2843,FA_out_2843}=REGS_58+REGS_121+REGS_188;
  assign {FA_cout_2844,FA_out_2844}=REGS_59+REGS_122+REGS_189;
  assign {FA_cout_2845,FA_out_2845}=REGS_60+REGS_123+REGS_190;
  assign {FA_cout_2846,FA_out_2846}=REGS_61+REGS_124+REGS_191;
  assign {FA_cout_2847,FA_out_2847}=REGS_62+REGS_125+REGS_192;
  assign {FA_cout_2848,FA_out_2848}=REGS_63+REGS_126+REGS_193;
  assign {FA_cout_2849,FA_out_2849}=REGS_64+REGS_127+REGS_194;
  assign {FA_cout_2850,FA_out_2850}=REGS_65+REGS_128+REGS_195;
  assign {FA_cout_2851,FA_out_2851}=REGS_66+REGS_129+REGS_196;
  assign {FA_cout_2852,FA_out_2852}=REGS_130+REGS_131+REGS_256;
  assign {FA_cout_2853,FA_out_2853}=REGS_132+REGS_133+REGS_260;
  assign {FA_cout_2854,FA_out_2854}=REGS_134+REGS_135+REGS_264;
  assign {FA_cout_2855,FA_out_2855}=REGS_136+REGS_197+REGS_268;
  assign {FA_cout_2856,FA_out_2856}=REGS_198+REGS_257+REGS_272;
  assign {FA_cout_2857,FA_out_2857}=REGS_206+REGS_286+REGS_340;
  assign {FA_cout_2858,FA_out_2858}=REGS_207+REGS_287+REGS_341;
  assign {FA_cout_2859,FA_out_2859}=REGS_208+REGS_288+REGS_342;
  assign {FA_cout_2860,FA_out_2860}=REGS_209+REGS_289+REGS_343;
  assign {FA_cout_2861,FA_out_2861}=REGS_210+REGS_290+REGS_344;
  assign {FA_cout_2862,FA_out_2862}=REGS_211+REGS_291+REGS_345;
  assign {FA_cout_2863,FA_out_2863}=REGS_212+REGS_292+REGS_346;
  assign {FA_cout_2864,FA_out_2864}=REGS_213+REGS_293+REGS_347;
  assign {FA_cout_2865,FA_out_2865}=REGS_214+REGS_294+REGS_348;
  assign {FA_cout_2866,FA_out_2866}=REGS_215+REGS_295+REGS_349;
  assign {FA_cout_2867,FA_out_2867}=REGS_216+REGS_296+REGS_350;
  assign {FA_cout_2868,FA_out_2868}=REGS_217+REGS_297+REGS_351;
  assign {FA_cout_2869,FA_out_2869}=REGS_218+REGS_298+REGS_352;
  assign {FA_cout_2870,FA_out_2870}=REGS_219+REGS_299+REGS_353;
  assign {FA_cout_2871,FA_out_2871}=REGS_220+REGS_300+REGS_354;
  assign {FA_cout_2872,FA_out_2872}=REGS_221+REGS_301+REGS_355;
  assign {FA_cout_2873,FA_out_2873}=REGS_222+REGS_302+REGS_356;
  assign {FA_cout_2874,FA_out_2874}=REGS_223+REGS_303+REGS_357;
  assign {FA_cout_2875,FA_out_2875}=REGS_224+REGS_304+REGS_358;
  assign {FA_cout_2876,FA_out_2876}=REGS_225+REGS_305+REGS_359;
  assign {FA_cout_2877,FA_out_2877}=REGS_226+REGS_306+REGS_360;
  assign {FA_cout_2878,FA_out_2878}=REGS_227+REGS_307+REGS_361;
  assign {FA_cout_2879,FA_out_2879}=REGS_228+REGS_308+REGS_362;
  assign {FA_cout_2880,FA_out_2880}=REGS_229+REGS_309+REGS_363;
  assign {FA_cout_2881,FA_out_2881}=REGS_230+REGS_310+REGS_364;
  assign {FA_cout_2882,FA_out_2882}=REGS_231+REGS_311+REGS_365;
  assign {FA_cout_2883,FA_out_2883}=REGS_232+REGS_312+REGS_366;
  assign {FA_cout_2884,FA_out_2884}=REGS_233+REGS_313+REGS_367;
  assign {FA_cout_2885,FA_out_2885}=REGS_234+REGS_314+REGS_368;
  assign {FA_cout_2886,FA_out_2886}=REGS_235+REGS_315+REGS_369;
  assign {FA_cout_2887,FA_out_2887}=REGS_236+REGS_316+REGS_370;
  assign {FA_cout_2888,FA_out_2888}=REGS_237+REGS_317+REGS_371;
  assign {FA_cout_2889,FA_out_2889}=REGS_238+REGS_318+REGS_372;
  assign {FA_cout_2890,FA_out_2890}=REGS_239+REGS_319+REGS_373;
  assign {FA_cout_2891,FA_out_2891}=REGS_240+REGS_320+REGS_374;
  assign {FA_cout_2892,FA_out_2892}=REGS_241+REGS_321+REGS_375;
  assign {FA_cout_2893,FA_out_2893}=REGS_242+REGS_322+REGS_376;
  assign {FA_cout_2894,FA_out_2894}=REGS_243+REGS_323+REGS_377;
  assign {FA_cout_2895,FA_out_2895}=REGS_244+REGS_324+REGS_378;
  assign {FA_cout_2896,FA_out_2896}=REGS_245+REGS_325+REGS_379;
  assign {FA_cout_2897,FA_out_2897}=REGS_246+REGS_326+REGS_380;
  assign {FA_cout_2898,FA_out_2898}=REGS_247+REGS_327+REGS_381;
  assign {FA_cout_2899,FA_out_2899}=REGS_248+REGS_328+REGS_382;
  assign {FA_cout_2900,FA_out_2900}=REGS_249+REGS_329+REGS_383;
  assign {FA_cout_2901,FA_out_2901}=REGS_250+REGS_330+REGS_384;
  assign {FA_cout_2902,FA_out_2902}=REGS_251+REGS_331+REGS_385;
  assign {FA_cout_2903,FA_out_2903}=REGS_252+REGS_332+REGS_386;
  assign {FA_cout_2904,FA_out_2904}=REGS_253+REGS_333+REGS_387;
  assign {FA_cout_2905,FA_out_2905}=REGS_254+REGS_334+REGS_388;
  assign {FA_cout_2906,FA_out_2906}=REGS_255+REGS_335+REGS_389;
  assign {FA_cout_2907,FA_out_2907}=REGS_258+REGS_261+REGS_276;
  assign {FA_cout_2908,FA_out_2908}=REGS_259+REGS_390+REGS_395;
  assign {FA_cout_2909,FA_out_2909}=REGS_262+REGS_265+REGS_280;
  assign {FA_cout_2910,FA_out_2910}=REGS_263+REGS_396+REGS_401;
  assign {FA_cout_2911,FA_out_2911}=REGS_266+REGS_269+REGS_337;
  assign {FA_cout_2912,FA_out_2912}=REGS_267+REGS_402+REGS_407;
  assign {FA_cout_2913,FA_out_2913}=REGS_270+REGS_273+REGS_392;
  assign {FA_cout_2914,FA_out_2914}=REGS_271+REGS_408+REGS_413;
  assign {FA_cout_2915,FA_out_2915}=REGS_274+REGS_277+REGS_398;
  assign {FA_cout_2916,FA_out_2916}=REGS_275+REGS_414+REGS_465;
  assign {FA_cout_2917,FA_out_2917}=REGS_278+REGS_281+REGS_404;
  assign {FA_cout_2918,FA_out_2918}=REGS_279+REGS_466+REGS_515;
  assign {FA_cout_2919,FA_out_2919}=REGS_282+REGS_338+REGS_410;
  assign {FA_cout_2920,FA_out_2920}=REGS_336+REGS_516+REGS_523;
  assign {FA_cout_2921,FA_out_2921}=REGS_339+REGS_393+REGS_416;
  assign {FA_cout_2922,FA_out_2922}=REGS_391+REGS_524+REGS_531;
  assign {FA_cout_2923,FA_out_2923}=REGS_394+REGS_399+REGS_468;
  assign {FA_cout_2924,FA_out_2924}=REGS_397+REGS_532+REGS_539;
  assign {FA_cout_2925,FA_out_2925}=REGS_400+REGS_405+REGS_518;
  assign {FA_cout_2926,FA_out_2926}=REGS_403+REGS_540+REGS_547;
  assign {FA_cout_2927,FA_out_2927}=REGS_406+REGS_411+REGS_526;
  assign {FA_cout_2928,FA_out_2928}=REGS_409+REGS_548+REGS_555;
  assign {FA_cout_2929,FA_out_2929}=REGS_412+REGS_417+REGS_534;
  assign {FA_cout_2930,FA_out_2930}=REGS_415+REGS_556+REGS_563;
  assign {FA_cout_2931,FA_out_2931}=REGS_418+REGS_469+REGS_542;
  assign {FA_cout_2932,FA_out_2932}=REGS_425+REGS_474+REGS_569;
  assign {FA_cout_2933,FA_out_2933}=REGS_426+REGS_475+REGS_570;
  assign {FA_cout_2934,FA_out_2934}=REGS_427+REGS_476+REGS_571;
  assign {FA_cout_2935,FA_out_2935}=REGS_428+REGS_477+REGS_572;
  assign {FA_cout_2936,FA_out_2936}=REGS_429+REGS_478+REGS_573;
  assign {FA_cout_2937,FA_out_2937}=REGS_430+REGS_479+REGS_574;
  assign {FA_cout_2938,FA_out_2938}=REGS_431+REGS_480+REGS_575;
  assign {FA_cout_2939,FA_out_2939}=REGS_432+REGS_481+REGS_576;
  assign {FA_cout_2940,FA_out_2940}=REGS_433+REGS_482+REGS_577;
  assign {FA_cout_2941,FA_out_2941}=REGS_434+REGS_483+REGS_578;
  assign {FA_cout_2942,FA_out_2942}=REGS_435+REGS_484+REGS_579;
  assign {FA_cout_2943,FA_out_2943}=REGS_436+REGS_485+REGS_580;
  assign {FA_cout_2944,FA_out_2944}=REGS_437+REGS_486+REGS_581;
  assign {FA_cout_2945,FA_out_2945}=REGS_438+REGS_487+REGS_582;
  assign {FA_cout_2946,FA_out_2946}=REGS_439+REGS_488+REGS_583;
  assign {FA_cout_2947,FA_out_2947}=REGS_440+REGS_489+REGS_584;
  assign {FA_cout_2948,FA_out_2948}=REGS_441+REGS_490+REGS_585;
  assign {FA_cout_2949,FA_out_2949}=REGS_442+REGS_491+REGS_586;
  assign {FA_cout_2950,FA_out_2950}=REGS_443+REGS_492+REGS_587;
  assign {FA_cout_2951,FA_out_2951}=REGS_444+REGS_493+REGS_588;
  assign {FA_cout_2952,FA_out_2952}=REGS_445+REGS_494+REGS_589;
  assign {FA_cout_2953,FA_out_2953}=REGS_446+REGS_495+REGS_590;
  assign {FA_cout_2954,FA_out_2954}=REGS_447+REGS_496+REGS_591;
  assign {FA_cout_2955,FA_out_2955}=REGS_448+REGS_497+REGS_592;
  assign {FA_cout_2956,FA_out_2956}=REGS_449+REGS_498+REGS_593;
  assign {FA_cout_2957,FA_out_2957}=REGS_450+REGS_499+REGS_594;
  assign {FA_cout_2958,FA_out_2958}=REGS_451+REGS_500+REGS_595;
  assign {FA_cout_2959,FA_out_2959}=REGS_452+REGS_501+REGS_596;
  assign {FA_cout_2960,FA_out_2960}=REGS_453+REGS_502+REGS_597;
  assign {FA_cout_2961,FA_out_2961}=REGS_454+REGS_503+REGS_598;
  assign {FA_cout_2962,FA_out_2962}=REGS_455+REGS_504+REGS_599;
  assign {FA_cout_2963,FA_out_2963}=REGS_456+REGS_505+REGS_600;
  assign {FA_cout_2964,FA_out_2964}=REGS_457+REGS_506+REGS_601;
  assign {FA_cout_2965,FA_out_2965}=REGS_458+REGS_507+REGS_602;
  assign {FA_cout_2966,FA_out_2966}=REGS_459+REGS_508+REGS_603;
  assign {FA_cout_2967,FA_out_2967}=REGS_460+REGS_509+REGS_604;
  assign {FA_cout_2968,FA_out_2968}=REGS_461+REGS_510+REGS_605;
  assign {FA_cout_2969,FA_out_2969}=REGS_462+REGS_511+REGS_606;
  assign {FA_cout_2970,FA_out_2970}=REGS_463+REGS_512+REGS_607;
  assign {FA_cout_2971,FA_out_2971}=REGS_464+REGS_513+REGS_608;
  assign {FA_cout_2972,FA_out_2972}=REGS_467+REGS_564+REGS_611;
  assign {FA_cout_2973,FA_out_2973}=REGS_470+REGS_519+REGS_550;
  assign {FA_cout_2974,FA_out_2974}=REGS_514+REGS_521+REGS_653;
  assign {FA_cout_2975,FA_out_2975}=REGS_517+REGS_612+REGS_656;
  assign {FA_cout_2976,FA_out_2976}=REGS_520+REGS_527+REGS_558;
  assign {FA_cout_2977,FA_out_2977}=REGS_522+REGS_529+REGS_663;
  assign {FA_cout_2978,FA_out_2978}=REGS_525+REGS_657+REGS_666;
  assign {FA_cout_2979,FA_out_2979}=REGS_528+REGS_535+REGS_566;
  assign {FA_cout_2980,FA_out_2980}=REGS_530+REGS_537+REGS_673;
  assign {FA_cout_2981,FA_out_2981}=REGS_533+REGS_667+REGS_676;
  assign {FA_cout_2982,FA_out_2982}=REGS_536+REGS_543+REGS_614;
  assign {FA_cout_2983,FA_out_2983}=REGS_538+REGS_545+REGS_683;
  assign {FA_cout_2984,FA_out_2984}=REGS_541+REGS_677+REGS_686;
  assign {FA_cout_2985,FA_out_2985}=REGS_544+REGS_551+REGS_659;
  assign {FA_cout_2986,FA_out_2986}=REGS_546+REGS_553+REGS_726;
  assign {FA_cout_2987,FA_out_2987}=REGS_549+REGS_687+REGS_729;
  assign {FA_cout_2988,FA_out_2988}=REGS_552+REGS_559+REGS_669;
  assign {FA_cout_2989,FA_out_2989}=REGS_554+REGS_561+REGS_767;
  assign {FA_cout_2990,FA_out_2990}=REGS_557+REGS_730+REGS_770;
  assign {FA_cout_2991,FA_out_2991}=REGS_560+REGS_567+REGS_679;
  assign {FA_cout_2992,FA_out_2992}=REGS_562+REGS_609+REGS_779;
  assign {FA_cout_2993,FA_out_2993}=REGS_565+REGS_771+REGS_782;
  assign {FA_cout_2994,FA_out_2994}=REGS_568+REGS_615+REGS_689;
  assign {FA_cout_2995,FA_out_2995}=REGS_610+REGS_654+REGS_791;
  assign {FA_cout_2996,FA_out_2996}=REGS_613+REGS_783+REGS_794;
  assign {FA_cout_2997,FA_out_2997}=REGS_616+REGS_660+REGS_732;
  assign {FA_cout_2998,FA_out_2998}=REGS_623+REGS_695+REGS_735;
  assign {FA_cout_2999,FA_out_2999}=REGS_624+REGS_696+REGS_736;
  assign {FA_cout_3000,FA_out_3000}=REGS_625+REGS_697+REGS_737;
  assign {FA_cout_3001,FA_out_3001}=REGS_626+REGS_698+REGS_738;
  assign {FA_cout_3002,FA_out_3002}=REGS_627+REGS_699+REGS_739;
  assign {FA_cout_3003,FA_out_3003}=REGS_628+REGS_700+REGS_740;
  assign {FA_cout_3004,FA_out_3004}=REGS_629+REGS_701+REGS_741;
  assign {FA_cout_3005,FA_out_3005}=REGS_630+REGS_702+REGS_742;
  assign {FA_cout_3006,FA_out_3006}=REGS_631+REGS_703+REGS_743;
  assign {FA_cout_3007,FA_out_3007}=REGS_632+REGS_704+REGS_744;
  assign {FA_cout_3008,FA_out_3008}=REGS_633+REGS_705+REGS_745;
  assign {FA_cout_3009,FA_out_3009}=REGS_634+REGS_706+REGS_746;
  assign {FA_cout_3010,FA_out_3010}=REGS_635+REGS_707+REGS_747;
  assign {FA_cout_3011,FA_out_3011}=REGS_636+REGS_708+REGS_748;
  assign {FA_cout_3012,FA_out_3012}=REGS_637+REGS_709+REGS_749;
  assign {FA_cout_3013,FA_out_3013}=REGS_638+REGS_710+REGS_750;
  assign {FA_cout_3014,FA_out_3014}=REGS_639+REGS_711+REGS_751;
  assign {FA_cout_3015,FA_out_3015}=REGS_640+REGS_712+REGS_752;
  assign {FA_cout_3016,FA_out_3016}=REGS_641+REGS_713+REGS_753;
  assign {FA_cout_3017,FA_out_3017}=REGS_642+REGS_714+REGS_754;
  assign {FA_cout_3018,FA_out_3018}=REGS_643+REGS_715+REGS_755;
  assign {FA_cout_3019,FA_out_3019}=REGS_644+REGS_716+REGS_756;
  assign {FA_cout_3020,FA_out_3020}=REGS_645+REGS_717+REGS_757;
  assign {FA_cout_3021,FA_out_3021}=REGS_646+REGS_718+REGS_758;
  assign {FA_cout_3022,FA_out_3022}=REGS_647+REGS_719+REGS_759;
  assign {FA_cout_3023,FA_out_3023}=REGS_648+REGS_720+REGS_760;
  assign {FA_cout_3024,FA_out_3024}=REGS_649+REGS_721+REGS_761;
  assign {FA_cout_3025,FA_out_3025}=REGS_650+REGS_722+REGS_762;
  assign {FA_cout_3026,FA_out_3026}=REGS_651+REGS_723+REGS_763;
  assign {FA_cout_3027,FA_out_3027}=REGS_652+REGS_724+REGS_764;
  assign {FA_cout_3028,FA_out_3028}=REGS_655+REGS_664+REGS_803;
  assign {FA_cout_3029,FA_out_3029}=REGS_658+REGS_795+REGS_806;
  assign {FA_cout_3030,FA_out_3030}=REGS_661+REGS_670+REGS_773;
  assign {FA_cout_3031,FA_out_3031}=REGS_662+REGS_765+REGS_776;
  assign {FA_cout_3032,FA_out_3032}=REGS_665+REGS_674+REGS_815;
  assign {FA_cout_3033,FA_out_3033}=REGS_668+REGS_807+REGS_818;
  assign {FA_cout_3034,FA_out_3034}=REGS_671+REGS_680+REGS_785;
  assign {FA_cout_3035,FA_out_3035}=REGS_672+REGS_777+REGS_788;
  assign {FA_cout_3036,FA_out_3036}=REGS_675+REGS_684+REGS_827;
  assign {FA_cout_3037,FA_out_3037}=REGS_678+REGS_819+REGS_830;
  assign {FA_cout_3038,FA_out_3038}=REGS_681+REGS_690+REGS_797;
  assign {FA_cout_3039,FA_out_3039}=REGS_682+REGS_789+REGS_800;
  assign {FA_cout_3040,FA_out_3040}=REGS_685+REGS_727+REGS_839;
  assign {FA_cout_3041,FA_out_3041}=REGS_688+REGS_831+REGS_842;
  assign {FA_cout_3042,FA_out_3042}=REGS_691+REGS_733+REGS_809;
  assign {FA_cout_3043,FA_out_3043}=REGS_725+REGS_801+REGS_812;
  assign {FA_cout_3044,FA_out_3044}=REGS_728+REGS_768+REGS_877;
  assign {FA_cout_3045,FA_out_3045}=REGS_731+REGS_843+REGS_880;
  assign {FA_cout_3046,FA_out_3046}=REGS_734+REGS_774+REGS_821;
  assign {FA_cout_3047,FA_out_3047}=REGS_766+REGS_813+REGS_824;
  assign {FA_cout_3048,FA_out_3048}=REGS_769+REGS_780+REGS_913;
  assign {FA_cout_3049,FA_out_3049}=REGS_772+REGS_881+REGS_916;
  assign {FA_cout_3050,FA_out_3050}=REGS_775+REGS_786+REGS_833;
  assign {FA_cout_3051,FA_out_3051}=REGS_778+REGS_825+REGS_836;
  assign {FA_cout_3052,FA_out_3052}=REGS_781+REGS_792+REGS_927;
  assign {FA_cout_3053,FA_out_3053}=REGS_784+REGS_917+REGS_930;
  assign {FA_cout_3054,FA_out_3054}=REGS_787+REGS_798+REGS_845;
  assign {FA_cout_3055,FA_out_3055}=REGS_790+REGS_837+REGS_874;
  assign {FA_cout_3056,FA_out_3056}=REGS_793+REGS_804+REGS_941;
  assign {FA_cout_3057,FA_out_3057}=REGS_796+REGS_931+REGS_944;
  assign {FA_cout_3058,FA_out_3058}=REGS_799+REGS_810+REGS_883;
  assign {FA_cout_3059,FA_out_3059}=REGS_802+REGS_875+REGS_910;
  assign {FA_cout_3060,FA_out_3060}=REGS_805+REGS_816+REGS_955;
  assign {FA_cout_3061,FA_out_3061}=REGS_808+REGS_945+REGS_958;
  assign {FA_cout_3062,FA_out_3062}=REGS_811+REGS_822+REGS_919;
  assign {FA_cout_3063,FA_out_3063}=REGS_814+REGS_911+REGS_924;
  assign {FA_cout_3064,FA_out_3064}=REGS_817+REGS_828+REGS_969;
  assign {FA_cout_3065,FA_out_3065}=REGS_820+REGS_959+REGS_972;
  assign {FA_cout_3066,FA_out_3066}=REGS_823+REGS_834+REGS_933;
  assign {FA_cout_3067,FA_out_3067}=REGS_826+REGS_925+REGS_938;
  assign {FA_cout_3068,FA_out_3068}=REGS_829+REGS_840+REGS_1002;
  assign {FA_cout_3069,FA_out_3069}=REGS_832+REGS_973+REGS_1005;
  assign {FA_cout_3070,FA_out_3070}=REGS_835+REGS_846+REGS_947;
  assign {FA_cout_3071,FA_out_3071}=REGS_838+REGS_939+REGS_952;
  assign {FA_cout_3072,FA_out_3072}=REGS_841+REGS_878+REGS_1033;
  assign {FA_cout_3073,FA_out_3073}=REGS_844+REGS_1006+REGS_1036;
  assign {FA_cout_3074,FA_out_3074}=REGS_847+REGS_884+REGS_961;
  assign {FA_cout_3075,FA_out_3075}=REGS_855+REGS_890+REGS_978;
  assign {FA_cout_3076,FA_out_3076}=REGS_856+REGS_891+REGS_979;
  assign {FA_cout_3077,FA_out_3077}=REGS_857+REGS_892+REGS_980;
  assign {FA_cout_3078,FA_out_3078}=REGS_858+REGS_893+REGS_981;
  assign {FA_cout_3079,FA_out_3079}=REGS_859+REGS_894+REGS_982;
  assign {FA_cout_3080,FA_out_3080}=REGS_860+REGS_895+REGS_983;
  assign {FA_cout_3081,FA_out_3081}=REGS_861+REGS_896+REGS_984;
  assign {FA_cout_3082,FA_out_3082}=REGS_862+REGS_897+REGS_985;
  assign {FA_cout_3083,FA_out_3083}=REGS_863+REGS_898+REGS_986;
  assign {FA_cout_3084,FA_out_3084}=REGS_864+REGS_899+REGS_987;
  assign {FA_cout_3085,FA_out_3085}=REGS_865+REGS_900+REGS_988;
  assign {FA_cout_3086,FA_out_3086}=REGS_866+REGS_901+REGS_989;
  assign {FA_cout_3087,FA_out_3087}=REGS_867+REGS_902+REGS_990;
  assign {FA_cout_3088,FA_out_3088}=REGS_868+REGS_903+REGS_991;
  assign {FA_cout_3089,FA_out_3089}=REGS_869+REGS_904+REGS_992;
  assign {FA_cout_3090,FA_out_3090}=REGS_870+REGS_905+REGS_993;
  assign {FA_cout_3091,FA_out_3091}=REGS_871+REGS_906+REGS_994;
  assign {FA_cout_3092,FA_out_3092}=REGS_872+REGS_907+REGS_995;
  assign {FA_cout_3093,FA_out_3093}=REGS_873+REGS_908+REGS_996;
  assign {FA_cout_3094,FA_out_3094}=REGS_876+REGS_953+REGS_966;
  assign {FA_cout_3095,FA_out_3095}=REGS_879+REGS_914+REGS_1049;
  assign {FA_cout_3096,FA_out_3096}=REGS_882+REGS_1037+REGS_1052;
  assign {FA_cout_3097,FA_out_3097}=REGS_885+REGS_920+REGS_975;
  assign {FA_cout_3098,FA_out_3098}=REGS_909+REGS_922+REGS_1027;
  assign {FA_cout_3099,FA_out_3099}=REGS_912+REGS_967+REGS_999;
  assign {FA_cout_3100,FA_out_3100}=REGS_915+REGS_928+REGS_1065;
  assign {FA_cout_3101,FA_out_3101}=REGS_918+REGS_1053+REGS_1068;
  assign {FA_cout_3102,FA_out_3102}=REGS_921+REGS_934+REGS_1008;
  assign {FA_cout_3103,FA_out_3103}=REGS_923+REGS_936+REGS_1043;
  assign {FA_cout_3104,FA_out_3104}=REGS_926+REGS_1000+REGS_1030;
  assign {FA_cout_3105,FA_out_3105}=REGS_929+REGS_942+REGS_1081;
  assign {FA_cout_3106,FA_out_3106}=REGS_932+REGS_1069+REGS_1084;
  assign {FA_cout_3107,FA_out_3107}=REGS_935+REGS_948+REGS_1039;
  assign {FA_cout_3108,FA_out_3108}=REGS_937+REGS_950+REGS_1059;
  assign {FA_cout_3109,FA_out_3109}=REGS_940+REGS_1031+REGS_1046;
  assign {FA_cout_3110,FA_out_3110}=REGS_943+REGS_956+REGS_1097;
  assign {FA_cout_3111,FA_out_3111}=REGS_946+REGS_1085+REGS_1100;
  assign {FA_cout_3112,FA_out_3112}=REGS_949+REGS_962+REGS_1055;
  assign {FA_cout_3113,FA_out_3113}=REGS_951+REGS_964+REGS_1075;
  assign {FA_cout_3114,FA_out_3114}=REGS_954+REGS_1047+REGS_1062;
  assign {FA_cout_3115,FA_out_3115}=REGS_957+REGS_970+REGS_1113;
  assign {FA_cout_3116,FA_out_3116}=REGS_960+REGS_1101+REGS_1116;
  assign {FA_cout_3117,FA_out_3117}=REGS_963+REGS_976+REGS_1071;
  assign {FA_cout_3118,FA_out_3118}=REGS_965+REGS_997+REGS_1091;
  assign {FA_cout_3119,FA_out_3119}=REGS_968+REGS_1063+REGS_1078;
  assign {FA_cout_3120,FA_out_3120}=REGS_971+REGS_1003+REGS_1129;
  assign {FA_cout_3121,FA_out_3121}=REGS_974+REGS_1117+REGS_1132;
  assign {FA_cout_3122,FA_out_3122}=REGS_977+REGS_1009+REGS_1087;
  assign {FA_cout_3123,FA_out_3123}=REGS_998+REGS_1028+REGS_1107;
  assign {FA_cout_3124,FA_out_3124}=REGS_1001+REGS_1079+REGS_1094;
  assign {FA_cout_3125,FA_out_3125}=REGS_1004+REGS_1034+REGS_1158;
  assign {FA_cout_3126,FA_out_3126}=REGS_1007+REGS_1133+REGS_1161;
  assign {FA_cout_3127,FA_out_3127}=REGS_1010+REGS_1040+REGS_1103;
  assign {FA_cout_3128,FA_out_3128}=REGS_1018+REGS_1142+REGS_1167;
  assign {FA_cout_3129,FA_out_3129}=REGS_1019+REGS_1143+REGS_1168;
  assign {FA_cout_3130,FA_out_3130}=REGS_1020+REGS_1144+REGS_1169;
  assign {FA_cout_3131,FA_out_3131}=REGS_1021+REGS_1145+REGS_1170;
  assign {FA_cout_3132,FA_out_3132}=REGS_1022+REGS_1146+REGS_1171;
  assign {FA_cout_3133,FA_out_3133}=REGS_1023+REGS_1147+REGS_1172;
  assign {FA_cout_3134,FA_out_3134}=REGS_1024+REGS_1148+REGS_1173;
  assign {FA_cout_3135,FA_out_3135}=REGS_1025+REGS_1149+REGS_1174;
  assign {FA_cout_3136,FA_out_3136}=REGS_1026+REGS_1150+REGS_1175;
  assign {FA_cout_3137,FA_out_3137}=REGS_1029+REGS_1044+REGS_1123;
  assign {FA_cout_3138,FA_out_3138}=REGS_1032+REGS_1095+REGS_1110;
  assign {FA_cout_3139,FA_out_3139}=REGS_1035+REGS_1050+REGS_1184;
  assign {FA_cout_3140,FA_out_3140}=REGS_1038+REGS_1162+REGS_1187;
  assign {FA_cout_3141,FA_out_3141}=REGS_1041+REGS_1056+REGS_1119;
  assign {FA_cout_3142,FA_out_3142}=REGS_1042+REGS_1176+REGS_1193;
  assign {FA_cout_3143,FA_out_3143}=REGS_1045+REGS_1060+REGS_1152;
  assign {FA_cout_3144,FA_out_3144}=REGS_1048+REGS_1111+REGS_1126;
  assign {FA_cout_3145,FA_out_3145}=REGS_1051+REGS_1066+REGS_1202;
  assign {FA_cout_3146,FA_out_3146}=REGS_1054+REGS_1188+REGS_1205;
  assign {FA_cout_3147,FA_out_3147}=REGS_1057+REGS_1072+REGS_1135;
  assign {FA_cout_3148,FA_out_3148}=REGS_1058+REGS_1194+REGS_1211;
  assign {FA_cout_3149,FA_out_3149}=REGS_1061+REGS_1076+REGS_1178;
  assign {FA_cout_3150,FA_out_3150}=REGS_1064+REGS_1127+REGS_1155;
  assign {FA_cout_3151,FA_out_3151}=REGS_1067+REGS_1082+REGS_1220;
  assign {FA_cout_3152,FA_out_3152}=REGS_1070+REGS_1206+REGS_1223;
  assign {FA_cout_3153,FA_out_3153}=REGS_1073+REGS_1088+REGS_1164;
  assign {FA_cout_3154,FA_out_3154}=REGS_1074+REGS_1212+REGS_1229;
  assign {FA_cout_3155,FA_out_3155}=REGS_1077+REGS_1092+REGS_1196;
  assign {FA_cout_3156,FA_out_3156}=REGS_1080+REGS_1156+REGS_1181;
  assign {FA_cout_3157,FA_out_3157}=REGS_1083+REGS_1098+REGS_1238;
  assign {FA_cout_3158,FA_out_3158}=REGS_1086+REGS_1224+REGS_1241;
  assign {FA_cout_3159,FA_out_3159}=REGS_1089+REGS_1104+REGS_1190;
  assign {FA_cout_3160,FA_out_3160}=REGS_1090+REGS_1230+REGS_1252;
  assign {FA_cout_3161,FA_out_3161}=REGS_1093+REGS_1108+REGS_1214;
  assign {FA_cout_3162,FA_out_3162}=REGS_1096+REGS_1182+REGS_1199;
  assign {FA_cout_3163,FA_out_3163}=REGS_1099+REGS_1114+REGS_1260;
  assign {FA_cout_3164,FA_out_3164}=REGS_1102+REGS_1242+REGS_1263;
  assign {FA_cout_3165,FA_out_3165}=REGS_1105+REGS_1120+REGS_1208;
  assign {FA_cout_3166,FA_out_3166}=REGS_1106+REGS_1253+REGS_1270;
  assign {FA_cout_3167,FA_out_3167}=REGS_1109+REGS_1124+REGS_1232;
  assign {FA_cout_3168,FA_out_3168}=REGS_1112+REGS_1200+REGS_1217;
  assign {FA_cout_3169,FA_out_3169}=REGS_1115+REGS_1130+REGS_1277;
  assign {FA_cout_3170,FA_out_3170}=REGS_1118+REGS_1264+REGS_1279;
  assign {FA_cout_3171,FA_out_3171}=REGS_1121+REGS_1136+REGS_1226;
  assign {FA_cout_3172,FA_out_3172}=REGS_1122+REGS_1271+REGS_1285;
  assign {FA_cout_3173,FA_out_3173}=REGS_1125+REGS_1153+REGS_1255;
  assign {FA_cout_3174,FA_out_3174}=REGS_1128+REGS_1218+REGS_1235;
  assign {FA_cout_3175,FA_out_3175}=REGS_1131+REGS_1159+REGS_1290;
  assign {FA_cout_3176,FA_out_3176}=REGS_1134+REGS_1280+REGS_1300;
  assign {FA_cout_3177,FA_out_3177}=REGS_1137+REGS_1165+REGS_1244;
  assign {FA_cout_3178,FA_out_3178}=REGS_1151+REGS_1286+REGS_1295;
  assign {FA_cout_3179,FA_out_3179}=REGS_1154+REGS_1179+REGS_1287;
  assign {FA_cout_3180,FA_out_3180}=REGS_1157+REGS_1236+REGS_1258;
  assign {FA_cout_3181,FA_out_3181}=REGS_1166+REGS_1191+REGS_1281;
  assign {FA_cout_3182,FA_out_3182}=REGS_1180+REGS_1197+REGS_1296;
  assign {FA_cout_3183,FA_out_3183}=REGS_1192+REGS_1209+REGS_1292;
  assign {FA_cout_3184,FA_out_3184}=FA_cout_2794+FA_out_2795+REGS_199;
  assign {FA_cout_3185,FA_out_3185}=FA_cout_2795+FA_out_2796+REGS_200;
  assign {FA_cout_3186,FA_out_3186}=FA_cout_2796+FA_out_2797+REGS_201;
  assign {FA_cout_3187,FA_out_3187}=FA_cout_2797+FA_out_2798+REGS_202;
  assign {FA_cout_3188,FA_out_3188}=FA_cout_2798+FA_out_2799+HA_out_129;
  assign {FA_cout_3189,FA_out_3189}=FA_cout_2799+FA_out_2800+HA_cout_129;
  assign {FA_cout_3190,FA_out_3190}=FA_cout_2800+FA_out_2801+HA_cout_130;
  assign {FA_cout_3191,FA_out_3191}=FA_cout_2801+FA_out_2802+HA_cout_131;
  assign {FA_cout_3192,FA_out_3192}=FA_cout_2802+FA_out_2803+FA_cout_2857;
  assign {FA_cout_3193,FA_out_3193}=FA_cout_2803+FA_out_2804+FA_cout_2858;
  assign {FA_cout_3194,FA_out_3194}=FA_cout_2804+FA_out_2805+FA_cout_2859;
  assign {FA_cout_3195,FA_out_3195}=FA_cout_2805+FA_out_2806+FA_cout_2860;
  assign {FA_cout_3196,FA_out_3196}=FA_cout_2806+FA_out_2807+FA_cout_2861;
  assign {FA_cout_3197,FA_out_3197}=FA_cout_2807+FA_out_2808+FA_cout_2862;
  assign {FA_cout_3198,FA_out_3198}=FA_cout_2808+FA_out_2809+FA_cout_2863;
  assign {FA_cout_3199,FA_out_3199}=FA_cout_2809+FA_out_2810+FA_cout_2864;
  assign {FA_cout_3200,FA_out_3200}=FA_cout_2810+FA_out_2811+FA_cout_2865;
  assign {FA_cout_3201,FA_out_3201}=FA_cout_2811+FA_out_2812+FA_cout_2866;
  assign {FA_cout_3202,FA_out_3202}=FA_cout_2812+FA_out_2813+FA_cout_2867;
  assign {FA_cout_3203,FA_out_3203}=FA_cout_2813+FA_out_2814+FA_cout_2868;
  assign {FA_cout_3204,FA_out_3204}=FA_cout_2814+FA_out_2815+FA_cout_2869;
  assign {FA_cout_3205,FA_out_3205}=FA_cout_2815+FA_out_2816+FA_cout_2870;
  assign {FA_cout_3206,FA_out_3206}=FA_cout_2816+FA_out_2817+FA_cout_2871;
  assign {FA_cout_3207,FA_out_3207}=FA_cout_2817+FA_out_2818+FA_cout_2872;
  assign {FA_cout_3208,FA_out_3208}=FA_cout_2818+FA_out_2819+FA_cout_2873;
  assign {FA_cout_3209,FA_out_3209}=FA_cout_2819+FA_out_2820+FA_cout_2874;
  assign {FA_cout_3210,FA_out_3210}=FA_cout_2820+FA_out_2821+FA_cout_2875;
  assign {FA_cout_3211,FA_out_3211}=FA_cout_2821+FA_out_2822+FA_cout_2876;
  assign {FA_cout_3212,FA_out_3212}=FA_cout_2822+FA_out_2823+FA_cout_2877;
  assign {FA_cout_3213,FA_out_3213}=FA_cout_2823+FA_out_2824+FA_cout_2878;
  assign {FA_cout_3214,FA_out_3214}=FA_cout_2824+FA_out_2825+FA_cout_2879;
  assign {FA_cout_3215,FA_out_3215}=FA_cout_2825+FA_out_2826+FA_cout_2880;
  assign {FA_cout_3216,FA_out_3216}=FA_cout_2826+FA_out_2827+FA_cout_2881;
  assign {FA_cout_3217,FA_out_3217}=FA_cout_2827+FA_out_2828+FA_cout_2882;
  assign {FA_cout_3218,FA_out_3218}=FA_cout_2828+FA_out_2829+FA_cout_2883;
  assign {FA_cout_3219,FA_out_3219}=FA_cout_2829+FA_out_2830+FA_cout_2884;
  assign {FA_cout_3220,FA_out_3220}=FA_cout_2830+FA_out_2831+FA_cout_2885;
  assign {FA_cout_3221,FA_out_3221}=FA_cout_2831+FA_out_2832+FA_cout_2886;
  assign {FA_cout_3222,FA_out_3222}=FA_cout_2832+FA_out_2833+FA_cout_2887;
  assign {FA_cout_3223,FA_out_3223}=FA_cout_2833+FA_out_2834+FA_cout_2888;
  assign {FA_cout_3224,FA_out_3224}=FA_cout_2834+FA_out_2835+FA_cout_2889;
  assign {FA_cout_3225,FA_out_3225}=FA_cout_2835+FA_out_2836+FA_cout_2890;
  assign {FA_cout_3226,FA_out_3226}=FA_cout_2836+FA_out_2837+FA_cout_2891;
  assign {FA_cout_3227,FA_out_3227}=FA_cout_2837+FA_out_2838+FA_cout_2892;
  assign {FA_cout_3228,FA_out_3228}=FA_cout_2838+FA_out_2839+FA_cout_2893;
  assign {FA_cout_3229,FA_out_3229}=FA_cout_2839+FA_out_2840+FA_cout_2894;
  assign {FA_cout_3230,FA_out_3230}=FA_cout_2840+FA_out_2841+FA_cout_2895;
  assign {FA_cout_3231,FA_out_3231}=FA_cout_2841+FA_out_2842+FA_cout_2896;
  assign {FA_cout_3232,FA_out_3232}=FA_cout_2842+FA_out_2843+FA_cout_2897;
  assign {FA_cout_3233,FA_out_3233}=FA_cout_2843+FA_out_2844+FA_cout_2898;
  assign {FA_cout_3234,FA_out_3234}=FA_cout_2844+FA_out_2845+FA_cout_2899;
  assign {FA_cout_3235,FA_out_3235}=FA_cout_2845+FA_out_2846+FA_cout_2900;
  assign {FA_cout_3236,FA_out_3236}=FA_cout_2846+FA_out_2847+FA_cout_2901;
  assign {FA_cout_3237,FA_out_3237}=FA_cout_2847+FA_out_2848+FA_cout_2902;
  assign {FA_cout_3238,FA_out_3238}=FA_cout_2848+FA_out_2849+FA_cout_2903;
  assign {FA_cout_3239,FA_out_3239}=FA_cout_2849+FA_out_2850+FA_cout_2904;
  assign {FA_cout_3240,FA_out_3240}=FA_cout_2850+FA_out_2851+FA_cout_2905;
  assign {FA_cout_3241,FA_out_3241}=FA_cout_2851+FA_out_2852+FA_cout_2906;
  assign {FA_cout_3242,FA_out_3242}=FA_cout_2852+FA_out_2853+FA_cout_2908;
  assign {FA_cout_3243,FA_out_3243}=FA_cout_2853+FA_out_2854+FA_cout_2910;
  assign {FA_cout_3244,FA_out_3244}=FA_cout_2854+FA_out_2855+FA_cout_2912;
  assign {FA_cout_3245,FA_out_3245}=FA_cout_2855+FA_out_2856+FA_cout_2914;
  assign {FA_cout_3246,FA_out_3246}=FA_cout_2856+FA_out_2907+FA_cout_2916;
  assign {FA_cout_3247,FA_out_3247}=FA_cout_2907+FA_out_2909+FA_cout_2918;
  assign {FA_cout_3248,FA_out_3248}=FA_out_2865+HA_cout_132+HA_out_133;
  assign {FA_cout_3249,FA_out_3249}=FA_out_2866+HA_cout_133+HA_out_134;
  assign {FA_cout_3250,FA_out_3250}=FA_out_2867+HA_cout_134+FA_out_2932;
  assign {FA_cout_3251,FA_out_3251}=FA_out_2868+FA_cout_2932+FA_out_2933;
  assign {FA_cout_3252,FA_out_3252}=FA_out_2869+FA_cout_2933+FA_out_2934;
  assign {FA_cout_3253,FA_out_3253}=FA_out_2870+FA_cout_2934+FA_out_2935;
  assign {FA_cout_3254,FA_out_3254}=FA_out_2871+FA_cout_2935+FA_out_2936;
  assign {FA_cout_3255,FA_out_3255}=FA_out_2872+FA_cout_2936+FA_out_2937;
  assign {FA_cout_3256,FA_out_3256}=FA_out_2873+FA_cout_2937+FA_out_2938;
  assign {FA_cout_3257,FA_out_3257}=FA_out_2874+FA_cout_2938+FA_out_2939;
  assign {FA_cout_3258,FA_out_3258}=FA_out_2875+FA_cout_2939+FA_out_2940;
  assign {FA_cout_3259,FA_out_3259}=FA_out_2876+FA_cout_2940+FA_out_2941;
  assign {FA_cout_3260,FA_out_3260}=FA_out_2877+FA_cout_2941+FA_out_2942;
  assign {FA_cout_3261,FA_out_3261}=FA_out_2878+FA_cout_2942+FA_out_2943;
  assign {FA_cout_3262,FA_out_3262}=FA_out_2879+FA_cout_2943+FA_out_2944;
  assign {FA_cout_3263,FA_out_3263}=FA_out_2880+FA_cout_2944+FA_out_2945;
  assign {FA_cout_3264,FA_out_3264}=FA_out_2881+FA_cout_2945+FA_out_2946;
  assign {FA_cout_3265,FA_out_3265}=FA_out_2882+FA_cout_2946+FA_out_2947;
  assign {FA_cout_3266,FA_out_3266}=FA_out_2883+FA_cout_2947+FA_out_2948;
  assign {FA_cout_3267,FA_out_3267}=FA_out_2884+FA_cout_2948+FA_out_2949;
  assign {FA_cout_3268,FA_out_3268}=FA_out_2885+FA_cout_2949+FA_out_2950;
  assign {FA_cout_3269,FA_out_3269}=FA_out_2886+FA_cout_2950+FA_out_2951;
  assign {FA_cout_3270,FA_out_3270}=FA_out_2887+FA_cout_2951+FA_out_2952;
  assign {FA_cout_3271,FA_out_3271}=FA_out_2888+FA_cout_2952+FA_out_2953;
  assign {FA_cout_3272,FA_out_3272}=FA_out_2889+FA_cout_2953+FA_out_2954;
  assign {FA_cout_3273,FA_out_3273}=FA_out_2890+FA_cout_2954+FA_out_2955;
  assign {FA_cout_3274,FA_out_3274}=FA_out_2891+FA_cout_2955+FA_out_2956;
  assign {FA_cout_3275,FA_out_3275}=FA_out_2892+FA_cout_2956+FA_out_2957;
  assign {FA_cout_3276,FA_out_3276}=FA_out_2893+FA_cout_2957+FA_out_2958;
  assign {FA_cout_3277,FA_out_3277}=FA_out_2894+FA_cout_2958+FA_out_2959;
  assign {FA_cout_3278,FA_out_3278}=FA_out_2895+FA_cout_2959+FA_out_2960;
  assign {FA_cout_3279,FA_out_3279}=FA_out_2896+FA_cout_2960+FA_out_2961;
  assign {FA_cout_3280,FA_out_3280}=FA_out_2897+FA_cout_2961+FA_out_2962;
  assign {FA_cout_3281,FA_out_3281}=FA_out_2898+FA_cout_2962+FA_out_2963;
  assign {FA_cout_3282,FA_out_3282}=FA_out_2899+FA_cout_2963+FA_out_2964;
  assign {FA_cout_3283,FA_out_3283}=FA_out_2900+FA_cout_2964+FA_out_2965;
  assign {FA_cout_3284,FA_out_3284}=FA_out_2901+FA_cout_2965+FA_out_2966;
  assign {FA_cout_3285,FA_out_3285}=FA_out_2902+FA_cout_2966+FA_out_2967;
  assign {FA_cout_3286,FA_out_3286}=FA_out_2903+FA_cout_2967+FA_out_2968;
  assign {FA_cout_3287,FA_out_3287}=FA_out_2904+FA_cout_2968+FA_out_2969;
  assign {FA_cout_3288,FA_out_3288}=FA_out_2905+FA_cout_2969+FA_out_2970;
  assign {FA_cout_3289,FA_out_3289}=FA_out_2906+FA_cout_2970+FA_out_2971;
  assign {FA_cout_3290,FA_out_3290}=FA_out_2908+FA_cout_2971+FA_out_2974;
  assign {FA_cout_3291,FA_out_3291}=FA_cout_2909+FA_out_2911+FA_cout_2920;
  assign {FA_cout_3292,FA_out_3292}=FA_out_2910+FA_cout_2974+FA_out_2977;
  assign {FA_cout_3293,FA_out_3293}=FA_cout_2911+FA_out_2913+FA_cout_2922;
  assign {FA_cout_3294,FA_out_3294}=FA_out_2912+FA_cout_2977+FA_out_2980;
  assign {FA_cout_3295,FA_out_3295}=FA_cout_2913+FA_out_2915+FA_cout_2924;
  assign {FA_cout_3296,FA_out_3296}=FA_out_2914+FA_cout_2980+FA_out_2983;
  assign {FA_cout_3297,FA_out_3297}=FA_cout_2915+FA_out_2917+FA_cout_2926;
  assign {FA_cout_3298,FA_out_3298}=FA_out_2916+FA_cout_2983+FA_out_2986;
  assign {FA_cout_3299,FA_out_3299}=FA_cout_2917+FA_out_2919+FA_cout_2928;
  assign {FA_cout_3300,FA_out_3300}=FA_out_2918+FA_cout_2986+FA_out_2989;
  assign {FA_cout_3301,FA_out_3301}=FA_cout_2919+FA_out_2921+FA_cout_2930;
  assign {FA_cout_3302,FA_out_3302}=FA_out_2920+FA_cout_2989+FA_out_2992;
  assign {FA_cout_3303,FA_out_3303}=FA_cout_2921+FA_out_2923+FA_cout_2972;
  assign {FA_cout_3304,FA_out_3304}=FA_out_2922+FA_cout_2992+FA_out_2995;
  assign {FA_cout_3305,FA_out_3305}=FA_cout_2923+FA_out_2925+FA_cout_2975;
  assign {FA_cout_3306,FA_out_3306}=FA_out_2924+FA_cout_2995+FA_out_3028;
  assign {FA_cout_3307,FA_out_3307}=FA_cout_2925+FA_out_2927+FA_cout_2978;
  assign {FA_cout_3308,FA_out_3308}=FA_out_2926+FA_cout_3028+FA_out_3032;
  assign {FA_cout_3309,FA_out_3309}=FA_cout_2927+FA_out_2929+FA_cout_2981;
  assign {FA_cout_3310,FA_out_3310}=FA_out_2928+FA_cout_3032+FA_out_3036;
  assign {FA_cout_3311,FA_out_3311}=FA_cout_2929+FA_out_2931+FA_cout_2984;
  assign {FA_cout_3312,FA_out_3312}=FA_out_2930+FA_cout_3036+FA_out_3040;
  assign {FA_cout_3313,FA_out_3313}=FA_cout_2931+FA_out_2973+FA_cout_2987;
  assign {FA_cout_3314,FA_out_3314}=FA_out_2972+FA_cout_3040+FA_out_3044;
  assign {FA_cout_3315,FA_out_3315}=FA_cout_2973+FA_out_2976+FA_cout_2990;
  assign {FA_cout_3316,FA_out_3316}=FA_out_2975+FA_cout_3044+FA_out_3048;
  assign {FA_cout_3317,FA_out_3317}=FA_cout_2976+FA_out_2979+FA_cout_2993;
  assign {FA_cout_3318,FA_out_3318}=FA_out_2978+FA_cout_3048+FA_out_3052;
  assign {FA_cout_3319,FA_out_3319}=FA_cout_2979+FA_out_2982+FA_cout_2996;
  assign {FA_cout_3320,FA_out_3320}=FA_out_2981+FA_cout_3052+FA_out_3056;
  assign {FA_cout_3321,FA_out_3321}=FA_cout_2982+FA_out_2985+FA_cout_3029;
  assign {FA_cout_3322,FA_out_3322}=FA_out_2984+FA_cout_3056+FA_out_3060;
  assign {FA_cout_3323,FA_out_3323}=FA_cout_2985+FA_out_2988+FA_cout_3033;
  assign {FA_cout_3324,FA_out_3324}=FA_out_2987+FA_cout_3060+FA_out_3064;
  assign {FA_cout_3325,FA_out_3325}=FA_cout_2988+FA_out_2991+FA_cout_3037;
  assign {FA_cout_3326,FA_out_3326}=FA_out_2990+FA_cout_3064+FA_out_3068;
  assign {FA_cout_3327,FA_out_3327}=FA_cout_2991+FA_out_2994+FA_cout_3041;
  assign {FA_cout_3328,FA_out_3328}=FA_out_2993+FA_cout_3068+FA_out_3072;
  assign {FA_cout_3329,FA_out_3329}=FA_cout_2994+FA_out_2997+FA_cout_3045;
  assign {FA_cout_3330,FA_out_3330}=FA_out_2996+FA_cout_3072+FA_out_3095;
  assign {FA_cout_3331,FA_out_3331}=FA_cout_2997+FA_out_3030+FA_cout_3049;
  assign {FA_cout_3332,FA_out_3332}=FA_cout_3001+FA_out_3002+REGS_848;
  assign {FA_cout_3333,FA_out_3333}=FA_cout_3002+FA_out_3003+REGS_849;
  assign {FA_cout_3334,FA_out_3334}=FA_cout_3003+FA_out_3004+REGS_850;
  assign {FA_cout_3335,FA_out_3335}=FA_cout_3004+FA_out_3005+HA_out_138;
  assign {FA_cout_3336,FA_out_3336}=FA_cout_3005+FA_out_3006+HA_cout_138;
  assign {FA_cout_3337,FA_out_3337}=FA_cout_3006+FA_out_3007+HA_cout_139;
  assign {FA_cout_3338,FA_out_3338}=FA_cout_3007+FA_out_3008+HA_cout_140;
  assign {FA_cout_3339,FA_out_3339}=FA_cout_3008+FA_out_3009+HA_cout_141;
  assign {FA_cout_3340,FA_out_3340}=FA_cout_3009+FA_out_3010+FA_cout_3075;
  assign {FA_cout_3341,FA_out_3341}=FA_cout_3010+FA_out_3011+FA_cout_3076;
  assign {FA_cout_3342,FA_out_3342}=FA_cout_3011+FA_out_3012+FA_cout_3077;
  assign {FA_cout_3343,FA_out_3343}=FA_cout_3012+FA_out_3013+FA_cout_3078;
  assign {FA_cout_3344,FA_out_3344}=FA_cout_3013+FA_out_3014+FA_cout_3079;
  assign {FA_cout_3345,FA_out_3345}=FA_cout_3014+FA_out_3015+FA_cout_3080;
  assign {FA_cout_3346,FA_out_3346}=FA_cout_3015+FA_out_3016+FA_cout_3081;
  assign {FA_cout_3347,FA_out_3347}=FA_cout_3016+FA_out_3017+FA_cout_3082;
  assign {FA_cout_3348,FA_out_3348}=FA_cout_3017+FA_out_3018+FA_cout_3083;
  assign {FA_cout_3349,FA_out_3349}=FA_cout_3018+FA_out_3019+FA_cout_3084;
  assign {FA_cout_3350,FA_out_3350}=FA_cout_3019+FA_out_3020+FA_cout_3085;
  assign {FA_cout_3351,FA_out_3351}=FA_cout_3020+FA_out_3021+FA_cout_3086;
  assign {FA_cout_3352,FA_out_3352}=FA_cout_3021+FA_out_3022+FA_cout_3087;
  assign {FA_cout_3353,FA_out_3353}=FA_cout_3022+FA_out_3023+FA_cout_3088;
  assign {FA_cout_3354,FA_out_3354}=FA_cout_3023+FA_out_3024+FA_cout_3089;
  assign {FA_cout_3355,FA_out_3355}=FA_cout_3024+FA_out_3025+FA_cout_3090;
  assign {FA_cout_3356,FA_out_3356}=FA_cout_3025+FA_out_3026+FA_cout_3091;
  assign {FA_cout_3357,FA_out_3357}=FA_cout_3026+FA_out_3027+FA_cout_3092;
  assign {FA_cout_3358,FA_out_3358}=FA_cout_3027+FA_out_3031+FA_cout_3093;
  assign {FA_cout_3359,FA_out_3359}=FA_out_3029+FA_cout_3095+FA_out_3100;
  assign {FA_cout_3360,FA_out_3360}=FA_cout_3030+FA_out_3034+FA_cout_3053;
  assign {FA_cout_3361,FA_out_3361}=FA_cout_3031+FA_out_3035+FA_cout_3098;
  assign {FA_cout_3362,FA_out_3362}=FA_out_3033+FA_cout_3100+FA_out_3105;
  assign {FA_cout_3363,FA_out_3363}=FA_cout_3034+FA_out_3038+FA_cout_3057;
  assign {FA_cout_3364,FA_out_3364}=FA_cout_3035+FA_out_3039+FA_cout_3103;
  assign {FA_cout_3365,FA_out_3365}=FA_out_3037+FA_cout_3105+FA_out_3110;
  assign {FA_cout_3366,FA_out_3366}=FA_cout_3038+FA_out_3042+FA_cout_3061;
  assign {FA_cout_3367,FA_out_3367}=FA_cout_3039+FA_out_3043+FA_cout_3108;
  assign {FA_cout_3368,FA_out_3368}=FA_out_3041+FA_cout_3110+FA_out_3115;
  assign {FA_cout_3369,FA_out_3369}=FA_cout_3042+FA_out_3046+FA_cout_3065;
  assign {FA_cout_3370,FA_out_3370}=FA_cout_3043+FA_out_3047+FA_cout_3113;
  assign {FA_cout_3371,FA_out_3371}=FA_out_3045+FA_cout_3115+FA_out_3120;
  assign {FA_cout_3372,FA_out_3372}=FA_cout_3046+FA_out_3050+FA_cout_3069;
  assign {FA_cout_3373,FA_out_3373}=FA_cout_3047+FA_out_3051+FA_cout_3118;
  assign {FA_cout_3374,FA_out_3374}=FA_out_3049+FA_cout_3120+FA_out_3125;
  assign {FA_cout_3375,FA_out_3375}=FA_cout_3050+FA_out_3054+FA_cout_3073;
  assign {FA_cout_3376,FA_out_3376}=FA_cout_3051+FA_out_3055+FA_cout_3123;
  assign {FA_cout_3377,FA_out_3377}=FA_out_3053+FA_cout_3125+FA_out_3139;
  assign {FA_cout_3378,FA_out_3378}=FA_cout_3054+FA_out_3058+FA_cout_3096;
  assign {FA_cout_3379,FA_out_3379}=FA_cout_3055+FA_out_3059+FA_cout_3137;
  assign {FA_cout_3380,FA_out_3380}=FA_out_3057+FA_cout_3139+FA_out_3145;
  assign {FA_cout_3381,FA_out_3381}=FA_cout_3058+FA_out_3062+FA_cout_3101;
  assign {FA_cout_3382,FA_out_3382}=FA_cout_3059+FA_out_3063+FA_cout_3143;
  assign {FA_cout_3383,FA_out_3383}=FA_out_3061+FA_cout_3145+FA_out_3151;
  assign {FA_cout_3384,FA_out_3384}=FA_cout_3062+FA_out_3066+FA_cout_3106;
  assign {FA_cout_3385,FA_out_3385}=FA_cout_3063+FA_out_3067+FA_cout_3149;
  assign {FA_cout_3386,FA_out_3386}=FA_out_3065+FA_cout_3151+FA_out_3157;
  assign {FA_cout_3387,FA_out_3387}=FA_cout_3066+FA_out_3070+FA_cout_3111;
  assign {FA_cout_3388,FA_out_3388}=FA_cout_3067+FA_out_3071+FA_cout_3155;
  assign {FA_cout_3389,FA_out_3389}=FA_out_3069+FA_cout_3157+FA_out_3163;
  assign {FA_cout_3390,FA_out_3390}=FA_cout_3070+FA_out_3074+FA_cout_3116;
  assign {FA_cout_3391,FA_out_3391}=FA_cout_3071+FA_out_3094+FA_cout_3161;
  assign {FA_cout_3392,FA_out_3392}=FA_out_3073+FA_cout_3163+FA_out_3169;
  assign {FA_cout_3393,FA_out_3393}=FA_cout_3074+FA_out_3097+FA_cout_3121;
  assign {FA_cout_3394,FA_out_3394}=FA_cout_3094+FA_out_3099+FA_cout_3167;
  assign {FA_cout_3395,FA_out_3395}=FA_out_3096+FA_cout_3169+FA_out_3175;
  assign {FA_cout_3396,FA_out_3396}=FA_cout_3097+FA_out_3102+FA_cout_3126;
  assign {FA_cout_3397,FA_out_3397}=FA_out_3082+HA_cout_142+HA_out_143;
  assign {FA_cout_3398,FA_out_3398}=FA_out_3083+HA_cout_143+HA_out_144;
  assign {FA_cout_3399,FA_out_3399}=FA_out_3084+HA_cout_144+HA_out_145;
  assign {FA_cout_3400,FA_out_3400}=FA_out_3085+HA_cout_145+FA_out_3128;
  assign {FA_cout_3401,FA_out_3401}=FA_out_3086+FA_cout_3128+FA_out_3129;
  assign {FA_cout_3402,FA_out_3402}=FA_out_3087+FA_cout_3129+FA_out_3130;
  assign {FA_cout_3403,FA_out_3403}=FA_out_3088+FA_cout_3130+FA_out_3131;
  assign {FA_cout_3404,FA_out_3404}=FA_out_3089+FA_cout_3131+FA_out_3132;
  assign {FA_cout_3405,FA_out_3405}=FA_out_3090+FA_cout_3132+FA_out_3133;
  assign {FA_cout_3406,FA_out_3406}=FA_out_3091+FA_cout_3133+FA_out_3134;
  assign {FA_cout_3407,FA_out_3407}=FA_out_3092+FA_cout_3134+FA_out_3135;
  assign {FA_cout_3408,FA_out_3408}=FA_out_3093+FA_cout_3135+FA_out_3136;
  assign {FA_cout_3409,FA_out_3409}=FA_out_3098+FA_cout_3136+FA_out_3142;
  assign {FA_cout_3410,FA_out_3410}=FA_cout_3099+FA_out_3104+FA_cout_3173;
  assign {FA_cout_3411,FA_out_3411}=FA_out_3101+FA_cout_3175+HA_out_146;
  assign {FA_cout_3412,FA_out_3412}=FA_cout_3102+FA_out_3107+FA_cout_3140;
  assign {FA_cout_3413,FA_out_3413}=FA_out_3103+FA_cout_3142+FA_out_3148;
  assign {FA_cout_3414,FA_out_3414}=FA_cout_3104+FA_out_3109+FA_cout_3179;
  assign {FA_cout_3415,FA_out_3415}=FA_out_3106+HA_cout_146+HA_out_149;
  assign {FA_cout_3416,FA_out_3416}=FA_cout_3107+FA_out_3112+FA_cout_3146;
  assign {FA_cout_3417,FA_out_3417}=FA_out_3108+FA_cout_3148+FA_out_3154;
  assign {FA_cout_3418,FA_out_3418}=FA_cout_3109+FA_out_3114+FA_cout_3182;
  assign {FA_cout_3419,FA_out_3419}=FA_out_3111+HA_cout_149+HA_out_152;
  assign {FA_cout_3420,FA_out_3420}=FA_cout_3112+FA_out_3117+FA_cout_3152;
  assign {FA_cout_3421,FA_out_3421}=FA_out_3113+FA_cout_3154+FA_out_3160;
  assign {FA_cout_3422,FA_out_3422}=FA_cout_3114+FA_out_3119+HA_cout_150;
  assign {FA_cout_3423,FA_out_3423}=FA_out_3116+HA_cout_152+HA_out_155;
  assign {FA_cout_3424,FA_out_3424}=FA_cout_3117+FA_out_3122+FA_cout_3158;
  assign {FA_cout_3425,FA_out_3425}=FA_out_3118+FA_cout_3160+FA_out_3166;
  assign {FA_cout_3426,FA_out_3426}=FA_cout_3119+FA_out_3124+HA_cout_154;
  assign {FA_cout_3427,FA_out_3427}=FA_out_3121+HA_cout_155+HA_out_158;
  assign {FA_cout_3428,FA_out_3428}=FA_cout_3122+FA_out_3127+FA_cout_3164;
  assign {FA_cout_3429,FA_out_3429}=FA_out_3123+FA_cout_3166+FA_out_3172;
  assign {FA_cout_3430,FA_out_3430}=FA_cout_3124+FA_out_3138+HA_cout_157;
  assign {FA_cout_3431,FA_out_3431}=FA_out_3126+HA_cout_158+HA_out_162;
  assign {FA_cout_3432,FA_out_3432}=FA_cout_3127+FA_out_3141+FA_cout_3170;
  assign {FA_cout_3433,FA_out_3433}=FA_out_3137+FA_cout_3172+FA_out_3178;
  assign {FA_cout_3434,FA_out_3434}=FA_cout_3138+FA_out_3144+HA_cout_161;
  assign {FA_cout_3435,FA_out_3435}=FA_out_3140+HA_cout_162+REGS_1291;
  assign {FA_cout_3436,FA_out_3436}=FA_cout_3141+FA_out_3147+FA_cout_3176;
  assign {FA_cout_3437,FA_out_3437}=FA_out_3143+FA_cout_3178+REGS_1177;
  assign {FA_cout_3438,FA_out_3438}=FA_cout_3144+FA_out_3150+HA_cout_164;
  assign {FA_cout_3439,FA_out_3439}=FA_cout_3147+FA_out_3153+HA_cout_147;
  assign {FA_cout_3440,FA_out_3440}=FA_cout_3153+FA_out_3159+REGS_1207;
  assign {FA_cout_3441,FA_out_3441}=FA_cout_3159+FA_out_3165+REGS_1225;
  assign {FA_cout_3442,FA_out_3442}=FA_cout_3165+FA_out_3171+REGS_1243;
  assign {FA_cout_3443,FA_out_3443}=FA_cout_3171+FA_out_3177+REGS_1265;
  assign {FA_cout_3444,FA_out_3444}=FA_cout_3188+FA_out_3189+HA_out_130;
  assign {FA_cout_3445,FA_out_3445}=FA_cout_3189+FA_out_3190+HA_out_131;
  assign {FA_cout_3446,FA_out_3446}=FA_cout_3190+FA_out_3191+FA_out_2857;
  assign {FA_cout_3447,FA_out_3447}=FA_cout_3191+FA_out_3192+FA_out_2858;
  assign {FA_cout_3448,FA_out_3448}=FA_cout_3192+FA_out_3193+FA_out_2859;
  assign {FA_cout_3449,FA_out_3449}=FA_cout_3193+FA_out_3194+FA_out_2860;
  assign {FA_cout_3450,FA_out_3450}=FA_cout_3194+FA_out_3195+HA_out_172;
  assign {FA_cout_3451,FA_out_3451}=FA_cout_3195+FA_out_3196+HA_cout_172;
  assign {FA_cout_3452,FA_out_3452}=FA_cout_3196+FA_out_3197+HA_cout_173;
  assign {FA_cout_3453,FA_out_3453}=FA_cout_3197+FA_out_3198+HA_cout_174;
  assign {FA_cout_3454,FA_out_3454}=FA_cout_3198+FA_out_3199+HA_cout_175;
  assign {FA_cout_3455,FA_out_3455}=FA_cout_3199+FA_out_3200+FA_cout_3248;
  assign {FA_cout_3456,FA_out_3456}=FA_cout_3200+FA_out_3201+FA_cout_3249;
  assign {FA_cout_3457,FA_out_3457}=FA_cout_3201+FA_out_3202+FA_cout_3250;
  assign {FA_cout_3458,FA_out_3458}=FA_cout_3202+FA_out_3203+FA_cout_3251;
  assign {FA_cout_3459,FA_out_3459}=FA_cout_3203+FA_out_3204+FA_cout_3252;
  assign {FA_cout_3460,FA_out_3460}=FA_cout_3204+FA_out_3205+FA_cout_3253;
  assign {FA_cout_3461,FA_out_3461}=FA_cout_3205+FA_out_3206+FA_cout_3254;
  assign {FA_cout_3462,FA_out_3462}=FA_cout_3206+FA_out_3207+FA_cout_3255;
  assign {FA_cout_3463,FA_out_3463}=FA_cout_3207+FA_out_3208+FA_cout_3256;
  assign {FA_cout_3464,FA_out_3464}=FA_cout_3208+FA_out_3209+FA_cout_3257;
  assign {FA_cout_3465,FA_out_3465}=FA_cout_3209+FA_out_3210+FA_cout_3258;
  assign {FA_cout_3466,FA_out_3466}=FA_cout_3210+FA_out_3211+FA_cout_3259;
  assign {FA_cout_3467,FA_out_3467}=FA_cout_3211+FA_out_3212+FA_cout_3260;
  assign {FA_cout_3468,FA_out_3468}=FA_cout_3212+FA_out_3213+FA_cout_3261;
  assign {FA_cout_3469,FA_out_3469}=FA_cout_3213+FA_out_3214+FA_cout_3262;
  assign {FA_cout_3470,FA_out_3470}=FA_cout_3214+FA_out_3215+FA_cout_3263;
  assign {FA_cout_3471,FA_out_3471}=FA_cout_3215+FA_out_3216+FA_cout_3264;
  assign {FA_cout_3472,FA_out_3472}=FA_cout_3216+FA_out_3217+FA_cout_3265;
  assign {FA_cout_3473,FA_out_3473}=FA_cout_3217+FA_out_3218+FA_cout_3266;
  assign {FA_cout_3474,FA_out_3474}=FA_cout_3218+FA_out_3219+FA_cout_3267;
  assign {FA_cout_3475,FA_out_3475}=FA_cout_3219+FA_out_3220+FA_cout_3268;
  assign {FA_cout_3476,FA_out_3476}=FA_cout_3220+FA_out_3221+FA_cout_3269;
  assign {FA_cout_3477,FA_out_3477}=FA_cout_3221+FA_out_3222+FA_cout_3270;
  assign {FA_cout_3478,FA_out_3478}=FA_cout_3222+FA_out_3223+FA_cout_3271;
  assign {FA_cout_3479,FA_out_3479}=FA_cout_3223+FA_out_3224+FA_cout_3272;
  assign {FA_cout_3480,FA_out_3480}=FA_cout_3224+FA_out_3225+FA_cout_3273;
  assign {FA_cout_3481,FA_out_3481}=FA_cout_3225+FA_out_3226+FA_cout_3274;
  assign {FA_cout_3482,FA_out_3482}=FA_cout_3226+FA_out_3227+FA_cout_3275;
  assign {FA_cout_3483,FA_out_3483}=FA_cout_3227+FA_out_3228+FA_cout_3276;
  assign {FA_cout_3484,FA_out_3484}=FA_cout_3228+FA_out_3229+FA_cout_3277;
  assign {FA_cout_3485,FA_out_3485}=FA_cout_3229+FA_out_3230+FA_cout_3278;
  assign {FA_cout_3486,FA_out_3486}=FA_cout_3230+FA_out_3231+FA_cout_3279;
  assign {FA_cout_3487,FA_out_3487}=FA_cout_3231+FA_out_3232+FA_cout_3280;
  assign {FA_cout_3488,FA_out_3488}=FA_cout_3232+FA_out_3233+FA_cout_3281;
  assign {FA_cout_3489,FA_out_3489}=FA_cout_3233+FA_out_3234+FA_cout_3282;
  assign {FA_cout_3490,FA_out_3490}=FA_cout_3234+FA_out_3235+FA_cout_3283;
  assign {FA_cout_3491,FA_out_3491}=FA_cout_3235+FA_out_3236+FA_cout_3284;
  assign {FA_cout_3492,FA_out_3492}=FA_cout_3236+FA_out_3237+FA_cout_3285;
  assign {FA_cout_3493,FA_out_3493}=FA_cout_3237+FA_out_3238+FA_cout_3286;
  assign {FA_cout_3494,FA_out_3494}=FA_cout_3238+FA_out_3239+FA_cout_3287;
  assign {FA_cout_3495,FA_out_3495}=FA_cout_3239+FA_out_3240+FA_cout_3288;
  assign {FA_cout_3496,FA_out_3496}=FA_cout_3240+FA_out_3241+FA_cout_3289;
  assign {FA_cout_3497,FA_out_3497}=FA_cout_3241+FA_out_3242+FA_cout_3290;
  assign {FA_cout_3498,FA_out_3498}=FA_cout_3242+FA_out_3243+FA_cout_3292;
  assign {FA_cout_3499,FA_out_3499}=FA_cout_3243+FA_out_3244+FA_cout_3294;
  assign {FA_cout_3500,FA_out_3500}=FA_cout_3244+FA_out_3245+FA_cout_3296;
  assign {FA_cout_3501,FA_out_3501}=FA_cout_3245+FA_out_3246+FA_cout_3298;
  assign {FA_cout_3502,FA_out_3502}=FA_cout_3246+FA_out_3247+FA_cout_3300;
  assign {FA_cout_3503,FA_out_3503}=FA_cout_3247+FA_out_3291+FA_cout_3302;
  assign {FA_cout_3504,FA_out_3504}=FA_cout_3291+FA_out_3293+FA_cout_3304;
  assign {FA_cout_3505,FA_out_3505}=FA_out_3259+HA_cout_176+HA_out_177;
  assign {FA_cout_3506,FA_out_3506}=FA_out_3260+HA_cout_177+HA_out_178;
  assign {FA_cout_3507,FA_out_3507}=FA_out_3261+HA_cout_178+HA_out_179;
  assign {FA_cout_3508,FA_out_3508}=FA_out_3262+HA_cout_179+HA_out_180;
  assign {FA_cout_3509,FA_out_3509}=FA_out_3263+HA_cout_180+HA_out_181;
  assign {FA_cout_3510,FA_out_3510}=FA_out_3264+HA_cout_181+FA_out_3332;
  assign {FA_cout_3511,FA_out_3511}=FA_out_3265+FA_cout_3332+FA_out_3333;
  assign {FA_cout_3512,FA_out_3512}=FA_out_3266+FA_cout_3333+FA_out_3334;
  assign {FA_cout_3513,FA_out_3513}=FA_out_3267+FA_cout_3334+FA_out_3335;
  assign {FA_cout_3514,FA_out_3514}=FA_out_3268+FA_cout_3335+FA_out_3336;
  assign {FA_cout_3515,FA_out_3515}=FA_out_3269+FA_cout_3336+FA_out_3337;
  assign {FA_cout_3516,FA_out_3516}=FA_out_3270+FA_cout_3337+FA_out_3338;
  assign {FA_cout_3517,FA_out_3517}=FA_out_3271+FA_cout_3338+FA_out_3339;
  assign {FA_cout_3518,FA_out_3518}=FA_out_3272+FA_cout_3339+FA_out_3340;
  assign {FA_cout_3519,FA_out_3519}=FA_out_3273+FA_cout_3340+FA_out_3341;
  assign {FA_cout_3520,FA_out_3520}=FA_out_3274+FA_cout_3341+FA_out_3342;
  assign {FA_cout_3521,FA_out_3521}=FA_out_3275+FA_cout_3342+FA_out_3343;
  assign {FA_cout_3522,FA_out_3522}=FA_out_3276+FA_cout_3343+FA_out_3344;
  assign {FA_cout_3523,FA_out_3523}=FA_out_3277+FA_cout_3344+FA_out_3345;
  assign {FA_cout_3524,FA_out_3524}=FA_out_3278+FA_cout_3345+FA_out_3346;
  assign {FA_cout_3525,FA_out_3525}=FA_out_3279+FA_cout_3346+FA_out_3347;
  assign {FA_cout_3526,FA_out_3526}=FA_out_3280+FA_cout_3347+FA_out_3348;
  assign {FA_cout_3527,FA_out_3527}=FA_out_3281+FA_cout_3348+FA_out_3349;
  assign {FA_cout_3528,FA_out_3528}=FA_out_3282+FA_cout_3349+FA_out_3350;
  assign {FA_cout_3529,FA_out_3529}=FA_out_3283+FA_cout_3350+FA_out_3351;
  assign {FA_cout_3530,FA_out_3530}=FA_out_3284+FA_cout_3351+FA_out_3352;
  assign {FA_cout_3531,FA_out_3531}=FA_out_3285+FA_cout_3352+FA_out_3353;
  assign {FA_cout_3532,FA_out_3532}=FA_out_3286+FA_cout_3353+FA_out_3354;
  assign {FA_cout_3533,FA_out_3533}=FA_out_3287+FA_cout_3354+FA_out_3355;
  assign {FA_cout_3534,FA_out_3534}=FA_out_3288+FA_cout_3355+FA_out_3356;
  assign {FA_cout_3535,FA_out_3535}=FA_out_3289+FA_cout_3356+FA_out_3357;
  assign {FA_cout_3536,FA_out_3536}=FA_out_3290+FA_cout_3357+FA_out_3358;
  assign {FA_cout_3537,FA_out_3537}=FA_out_3292+FA_cout_3358+FA_out_3361;
  assign {FA_cout_3538,FA_out_3538}=FA_cout_3293+FA_out_3295+FA_cout_3306;
  assign {FA_cout_3539,FA_out_3539}=FA_out_3294+FA_cout_3361+FA_out_3364;
  assign {FA_cout_3540,FA_out_3540}=FA_cout_3295+FA_out_3297+FA_cout_3308;
  assign {FA_cout_3541,FA_out_3541}=FA_out_3296+FA_cout_3364+FA_out_3367;
  assign {FA_cout_3542,FA_out_3542}=FA_cout_3297+FA_out_3299+FA_cout_3310;
  assign {FA_cout_3543,FA_out_3543}=FA_out_3298+FA_cout_3367+FA_out_3370;
  assign {FA_cout_3544,FA_out_3544}=FA_cout_3299+FA_out_3301+FA_cout_3312;
  assign {FA_cout_3545,FA_out_3545}=FA_out_3300+FA_cout_3370+FA_out_3373;
  assign {FA_cout_3546,FA_out_3546}=FA_cout_3301+FA_out_3303+FA_cout_3314;
  assign {FA_cout_3547,FA_out_3547}=FA_out_3302+FA_cout_3373+FA_out_3376;
  assign {FA_cout_3548,FA_out_3548}=FA_cout_3303+FA_out_3305+FA_cout_3316;
  assign {FA_cout_3549,FA_out_3549}=FA_out_3304+FA_cout_3376+FA_out_3379;
  assign {FA_cout_3550,FA_out_3550}=FA_cout_3305+FA_out_3307+FA_cout_3318;
  assign {FA_cout_3551,FA_out_3551}=FA_out_3306+FA_cout_3379+FA_out_3382;
  assign {FA_cout_3552,FA_out_3552}=FA_cout_3307+FA_out_3309+FA_cout_3320;
  assign {FA_cout_3553,FA_out_3553}=FA_out_3308+FA_cout_3382+FA_out_3385;
  assign {FA_cout_3554,FA_out_3554}=FA_cout_3309+FA_out_3311+FA_cout_3322;
  assign {FA_cout_3555,FA_out_3555}=FA_out_3310+FA_cout_3385+FA_out_3388;
  assign {FA_cout_3556,FA_out_3556}=FA_cout_3311+FA_out_3313+FA_cout_3324;
  assign {FA_cout_3557,FA_out_3557}=FA_out_3312+FA_cout_3388+FA_out_3391;
  assign {FA_cout_3558,FA_out_3558}=FA_cout_3313+FA_out_3315+FA_cout_3326;
  assign {FA_cout_3559,FA_out_3559}=FA_out_3314+FA_cout_3391+FA_out_3394;
  assign {FA_cout_3560,FA_out_3560}=FA_cout_3315+FA_out_3317+FA_cout_3328;
  assign {FA_cout_3561,FA_out_3561}=FA_out_3316+FA_cout_3394+FA_out_3410;
  assign {FA_cout_3562,FA_out_3562}=FA_cout_3317+FA_out_3319+FA_cout_3330;
  assign {FA_cout_3563,FA_out_3563}=FA_out_3318+FA_cout_3410+FA_out_3414;
  assign {FA_cout_3564,FA_out_3564}=FA_cout_3319+FA_out_3321+FA_cout_3359;
  assign {FA_cout_3565,FA_out_3565}=FA_out_3320+FA_cout_3414+FA_out_3418;
  assign {FA_cout_3566,FA_out_3566}=FA_cout_3321+FA_out_3323+FA_cout_3362;
  assign {FA_cout_3567,FA_out_3567}=FA_out_3322+FA_cout_3418+FA_out_3422;
  assign {FA_cout_3568,FA_out_3568}=FA_cout_3323+FA_out_3325+FA_cout_3365;
  assign {FA_cout_3569,FA_out_3569}=FA_out_3324+FA_cout_3422+FA_out_3426;
  assign {FA_cout_3570,FA_out_3570}=FA_cout_3325+FA_out_3327+FA_cout_3368;
  assign {FA_cout_3571,FA_out_3571}=FA_out_3326+FA_cout_3426+FA_out_3430;
  assign {FA_cout_3572,FA_out_3572}=FA_cout_3327+FA_out_3329+FA_cout_3371;
  assign {FA_cout_3573,FA_out_3573}=FA_out_3328+FA_cout_3430+FA_out_3434;
  assign {FA_cout_3574,FA_out_3574}=FA_cout_3329+FA_out_3331+FA_cout_3374;
  assign {FA_cout_3575,FA_out_3575}=FA_out_3330+FA_cout_3434+FA_out_3438;
  assign {FA_cout_3576,FA_out_3576}=FA_cout_3331+FA_out_3360+FA_cout_3377;
  assign {FA_cout_3577,FA_out_3577}=FA_out_3359+FA_cout_3438+HA_out_188;
  assign {FA_cout_3578,FA_out_3578}=FA_cout_3360+FA_out_3363+FA_cout_3380;
  assign {FA_cout_3579,FA_out_3579}=FA_out_3362+HA_cout_188+HA_out_190;
  assign {FA_cout_3580,FA_out_3580}=FA_cout_3363+FA_out_3366+FA_cout_3383;
  assign {FA_cout_3581,FA_out_3581}=FA_out_3365+HA_cout_190+HA_out_192;
  assign {FA_cout_3582,FA_out_3582}=FA_cout_3366+FA_out_3369+FA_cout_3386;
  assign {FA_cout_3583,FA_out_3583}=FA_out_3368+HA_cout_192+HA_out_194;
  assign {FA_cout_3584,FA_out_3584}=FA_cout_3369+FA_out_3372+FA_cout_3389;
  assign {FA_cout_3585,FA_out_3585}=FA_out_3371+HA_cout_194+HA_out_196;
  assign {FA_cout_3586,FA_out_3586}=FA_cout_3372+FA_out_3375+FA_cout_3392;
  assign {FA_cout_3587,FA_out_3587}=FA_out_3374+HA_cout_196+HA_out_198;
  assign {FA_cout_3588,FA_out_3588}=FA_cout_3375+FA_out_3378+FA_cout_3395;
  assign {FA_cout_3589,FA_out_3589}=FA_out_3377+HA_cout_198+HA_out_200;
  assign {FA_cout_3590,FA_out_3590}=FA_cout_3378+FA_out_3381+FA_cout_3411;
  assign {FA_cout_3591,FA_out_3591}=FA_out_3380+HA_cout_200+HA_out_202;
  assign {FA_cout_3592,FA_out_3592}=FA_cout_3381+FA_out_3384+FA_cout_3415;
  assign {FA_cout_3593,FA_out_3593}=FA_out_3383+HA_cout_202+REGS_1237;
  assign {FA_cout_3594,FA_out_3594}=FA_cout_3384+FA_out_3387+FA_cout_3419;
  assign {FA_cout_3595,FA_out_3595}=FA_cout_3387+FA_out_3390+FA_cout_3423;
  assign {FA_cout_3596,FA_out_3596}=FA_cout_3390+FA_out_3393+FA_cout_3427;
  assign {FA_cout_3597,FA_out_3597}=FA_cout_3393+FA_out_3396+FA_cout_3431;
  assign {FA_cout_3598,FA_out_3598}=FA_cout_3396+FA_out_3412+FA_cout_3435;
  assign {FA_cout_3599,FA_out_3599}=FA_cout_3402+FA_out_3403+REGS_1247;
  assign {FA_cout_3600,FA_out_3600}=FA_cout_3403+FA_out_3404+REGS_1248;
  assign {FA_cout_3601,FA_out_3601}=FA_cout_3404+FA_out_3405+REGS_1249;
  assign {FA_cout_3602,FA_out_3602}=FA_cout_3405+FA_out_3406+HA_out_160;
  assign {FA_cout_3603,FA_out_3603}=FA_cout_3406+FA_out_3407+HA_out_206;
  assign {FA_cout_3604,FA_out_3604}=FA_cout_3407+FA_out_3408+HA_cout_206;
  assign {FA_cout_3605,FA_out_3605}=FA_cout_3408+FA_out_3409+REGS_1284;
  assign {FA_cout_3606,FA_out_3606}=FA_cout_3412+FA_out_3416+HA_cout_186;
  assign {FA_cout_3607,FA_out_3607}=FA_cout_3416+FA_out_3420+FA_out_3158;
  assign {FA_cout_3608,FA_out_3608}=FA_cout_3420+FA_out_3424+FA_out_3164;
  assign {FA_cout_3609,FA_out_3609}=FA_cout_3424+FA_out_3428+FA_out_3170;
  assign {FA_cout_3610,FA_out_3610}=FA_cout_3428+FA_out_3432+FA_out_3176;
  assign {FA_cout_3611,FA_out_3611}=FA_cout_3432+FA_out_3436+HA_out_147;
  assign {FA_cout_3612,FA_out_3612}=FA_cout_3436+FA_out_3439+REGS_1189;
  assign {FA_cout_3613,FA_out_3613}=FA_cout_3450+FA_out_3451+HA_out_173;
  assign {FA_cout_3614,FA_out_3614}=FA_cout_3451+FA_out_3452+HA_out_174;
  assign {FA_cout_3615,FA_out_3615}=FA_cout_3452+FA_out_3453+HA_out_175;
  assign {FA_cout_3616,FA_out_3616}=FA_cout_3453+FA_out_3454+FA_out_3248;
  assign {FA_cout_3617,FA_out_3617}=FA_cout_3454+FA_out_3455+FA_out_3249;
  assign {FA_cout_3618,FA_out_3618}=FA_cout_3455+FA_out_3456+FA_out_3250;
  assign {FA_cout_3619,FA_out_3619}=FA_cout_3456+FA_out_3457+FA_out_3251;
  assign {FA_cout_3620,FA_out_3620}=FA_cout_3457+FA_out_3458+FA_out_3252;
  assign {FA_cout_3621,FA_out_3621}=FA_cout_3458+FA_out_3459+FA_out_3253;
  assign {FA_cout_3622,FA_out_3622}=FA_cout_3459+FA_out_3460+HA_out_218;
  assign {FA_cout_3623,FA_out_3623}=FA_cout_3460+FA_out_3461+HA_cout_218;
  assign {FA_cout_3624,FA_out_3624}=FA_cout_3461+FA_out_3462+HA_cout_219;
  assign {FA_cout_3625,FA_out_3625}=FA_cout_3462+FA_out_3463+HA_cout_220;
  assign {FA_cout_3626,FA_out_3626}=FA_cout_3463+FA_out_3464+HA_cout_221;
  assign {FA_cout_3627,FA_out_3627}=FA_cout_3464+FA_out_3465+HA_cout_222;
  assign {FA_cout_3628,FA_out_3628}=FA_cout_3465+FA_out_3466+FA_cout_3505;
  assign {FA_cout_3629,FA_out_3629}=FA_cout_3466+FA_out_3467+FA_cout_3506;
  assign {FA_cout_3630,FA_out_3630}=FA_cout_3467+FA_out_3468+FA_cout_3507;
  assign {FA_cout_3631,FA_out_3631}=FA_cout_3468+FA_out_3469+FA_cout_3508;
  assign {FA_cout_3632,FA_out_3632}=FA_cout_3469+FA_out_3470+FA_cout_3509;
  assign {FA_cout_3633,FA_out_3633}=FA_cout_3470+FA_out_3471+FA_cout_3510;
  assign {FA_cout_3634,FA_out_3634}=FA_cout_3471+FA_out_3472+FA_cout_3511;
  assign {FA_cout_3635,FA_out_3635}=FA_cout_3472+FA_out_3473+FA_cout_3512;
  assign {FA_cout_3636,FA_out_3636}=FA_cout_3473+FA_out_3474+FA_cout_3513;
  assign {FA_cout_3637,FA_out_3637}=FA_cout_3474+FA_out_3475+FA_cout_3514;
  assign {FA_cout_3638,FA_out_3638}=FA_cout_3475+FA_out_3476+FA_cout_3515;
  assign {FA_cout_3639,FA_out_3639}=FA_cout_3476+FA_out_3477+FA_cout_3516;
  assign {FA_cout_3640,FA_out_3640}=FA_cout_3477+FA_out_3478+FA_cout_3517;
  assign {FA_cout_3641,FA_out_3641}=FA_cout_3478+FA_out_3479+FA_cout_3518;
  assign {FA_cout_3642,FA_out_3642}=FA_cout_3479+FA_out_3480+FA_cout_3519;
  assign {FA_cout_3643,FA_out_3643}=FA_cout_3480+FA_out_3481+FA_cout_3520;
  assign {FA_cout_3644,FA_out_3644}=FA_cout_3481+FA_out_3482+FA_cout_3521;
  assign {FA_cout_3645,FA_out_3645}=FA_cout_3482+FA_out_3483+FA_cout_3522;
  assign {FA_cout_3646,FA_out_3646}=FA_cout_3483+FA_out_3484+FA_cout_3523;
  assign {FA_cout_3647,FA_out_3647}=FA_cout_3484+FA_out_3485+FA_cout_3524;
  assign {FA_cout_3648,FA_out_3648}=FA_cout_3485+FA_out_3486+FA_cout_3525;
  assign {FA_cout_3649,FA_out_3649}=FA_cout_3486+FA_out_3487+FA_cout_3526;
  assign {FA_cout_3650,FA_out_3650}=FA_cout_3487+FA_out_3488+FA_cout_3527;
  assign {FA_cout_3651,FA_out_3651}=FA_cout_3488+FA_out_3489+FA_cout_3528;
  assign {FA_cout_3652,FA_out_3652}=FA_cout_3489+FA_out_3490+FA_cout_3529;
  assign {FA_cout_3653,FA_out_3653}=FA_cout_3490+FA_out_3491+FA_cout_3530;
  assign {FA_cout_3654,FA_out_3654}=FA_cout_3491+FA_out_3492+FA_cout_3531;
  assign {FA_cout_3655,FA_out_3655}=FA_cout_3492+FA_out_3493+FA_cout_3532;
  assign {FA_cout_3656,FA_out_3656}=FA_cout_3493+FA_out_3494+FA_cout_3533;
  assign {FA_cout_3657,FA_out_3657}=FA_cout_3494+FA_out_3495+FA_cout_3534;
  assign {FA_cout_3658,FA_out_3658}=FA_cout_3495+FA_out_3496+FA_cout_3535;
  assign {FA_cout_3659,FA_out_3659}=FA_cout_3496+FA_out_3497+FA_cout_3536;
  assign {FA_cout_3660,FA_out_3660}=FA_cout_3497+FA_out_3498+FA_cout_3537;
  assign {FA_cout_3661,FA_out_3661}=FA_cout_3498+FA_out_3499+FA_cout_3539;
  assign {FA_cout_3662,FA_out_3662}=FA_cout_3499+FA_out_3500+FA_cout_3541;
  assign {FA_cout_3663,FA_out_3663}=FA_cout_3500+FA_out_3501+FA_cout_3543;
  assign {FA_cout_3664,FA_out_3664}=FA_cout_3501+FA_out_3502+FA_cout_3545;
  assign {FA_cout_3665,FA_out_3665}=FA_cout_3502+FA_out_3503+FA_cout_3547;
  assign {FA_cout_3666,FA_out_3666}=FA_cout_3503+FA_out_3504+FA_cout_3549;
  assign {FA_cout_3667,FA_out_3667}=FA_cout_3504+FA_out_3538+FA_cout_3551;
  assign {FA_cout_3668,FA_out_3668}=FA_cout_3538+FA_out_3540+FA_cout_3553;
  assign {FA_cout_3669,FA_out_3669}=FA_out_3522+HA_cout_227+HA_out_228;
  assign {FA_cout_3670,FA_out_3670}=FA_out_3523+HA_cout_228+HA_out_229;
  assign {FA_cout_3671,FA_out_3671}=FA_out_3524+HA_cout_229+HA_out_230;
  assign {FA_cout_3672,FA_out_3672}=FA_out_3525+HA_cout_230+HA_out_231;
  assign {FA_cout_3673,FA_out_3673}=FA_out_3526+HA_cout_231+HA_out_232;
  assign {FA_cout_3674,FA_out_3674}=FA_out_3527+HA_cout_232+HA_out_233;
  assign {FA_cout_3675,FA_out_3675}=FA_out_3528+HA_cout_233+HA_out_234;
  assign {FA_cout_3676,FA_out_3676}=FA_out_3529+HA_cout_234+HA_out_235;
  assign {FA_cout_3677,FA_out_3677}=FA_out_3530+HA_cout_235+FA_out_3599;
  assign {FA_cout_3678,FA_out_3678}=FA_out_3531+FA_cout_3599+FA_out_3600;
  assign {FA_cout_3679,FA_out_3679}=FA_out_3532+FA_cout_3600+FA_out_3601;
  assign {FA_cout_3680,FA_out_3680}=FA_out_3533+FA_cout_3601+FA_out_3602;
  assign {FA_cout_3681,FA_out_3681}=FA_out_3534+FA_cout_3602+FA_out_3603;
  assign {FA_cout_3682,FA_out_3682}=FA_out_3535+FA_cout_3603+FA_out_3604;
  assign {FA_cout_3683,FA_out_3683}=FA_out_3536+FA_cout_3604+FA_out_3605;
  assign {FA_cout_3684,FA_out_3684}=FA_out_3537+FA_cout_3605+HA_out_236;
  assign {FA_cout_3685,FA_out_3685}=FA_out_3539+HA_cout_236+HA_out_237;
  assign {FA_cout_3686,FA_out_3686}=FA_cout_3540+FA_out_3542+FA_cout_3555;
  assign {FA_cout_3687,FA_out_3687}=FA_out_3541+HA_cout_237+HA_out_238;
  assign {FA_cout_3688,FA_out_3688}=FA_cout_3542+FA_out_3544+FA_cout_3557;
  assign {FA_cout_3689,FA_out_3689}=FA_out_3543+HA_cout_238+HA_out_239;
  assign {FA_cout_3690,FA_out_3690}=FA_cout_3544+FA_out_3546+FA_cout_3559;
  assign {FA_cout_3691,FA_out_3691}=FA_out_3545+HA_cout_239+HA_out_240;
  assign {FA_cout_3692,FA_out_3692}=FA_cout_3546+FA_out_3548+FA_cout_3561;
  assign {FA_cout_3693,FA_out_3693}=FA_out_3547+HA_cout_240+HA_out_241;
  assign {FA_cout_3694,FA_out_3694}=FA_cout_3548+FA_out_3550+FA_cout_3563;
  assign {FA_cout_3695,FA_out_3695}=FA_out_3549+HA_cout_241+HA_out_242;
  assign {FA_cout_3696,FA_out_3696}=FA_cout_3550+FA_out_3552+FA_cout_3565;
  assign {FA_cout_3697,FA_out_3697}=FA_out_3551+HA_cout_242+HA_out_243;
  assign {FA_cout_3698,FA_out_3698}=FA_cout_3552+FA_out_3554+FA_cout_3567;
  assign {FA_cout_3699,FA_out_3699}=FA_out_3553+HA_cout_243+HA_out_245;
  assign {FA_cout_3700,FA_out_3700}=FA_cout_3554+FA_out_3556+FA_cout_3569;
  assign {FA_cout_3701,FA_out_3701}=FA_out_3555+HA_cout_245+HA_out_247;
  assign {FA_cout_3702,FA_out_3702}=FA_cout_3556+FA_out_3558+FA_cout_3571;
  assign {FA_cout_3703,FA_out_3703}=FA_out_3557+HA_cout_247+HA_out_249;
  assign {FA_cout_3704,FA_out_3704}=FA_cout_3558+FA_out_3560+FA_cout_3573;
  assign {FA_cout_3705,FA_out_3705}=FA_out_3559+HA_cout_249+HA_out_251;
  assign {FA_cout_3706,FA_out_3706}=FA_cout_3560+FA_out_3562+FA_cout_3575;
  assign {FA_cout_3707,FA_out_3707}=FA_out_3561+HA_cout_251+HA_out_253;
  assign {FA_cout_3708,FA_out_3708}=FA_cout_3562+FA_out_3564+FA_cout_3577;
  assign {FA_cout_3709,FA_out_3709}=FA_out_3563+HA_cout_253+FA_out_3182;
  assign {FA_cout_3710,FA_out_3710}=FA_cout_3564+FA_out_3566+FA_cout_3579;
  assign {FA_cout_3711,FA_out_3711}=FA_cout_3566+FA_out_3568+FA_cout_3581;
  assign {FA_cout_3712,FA_out_3712}=FA_cout_3568+FA_out_3570+FA_cout_3583;
  assign {FA_cout_3713,FA_out_3713}=FA_cout_3570+FA_out_3572+FA_cout_3585;
  assign {FA_cout_3714,FA_out_3714}=FA_cout_3572+FA_out_3574+FA_cout_3587;
  assign {FA_cout_3715,FA_out_3715}=FA_cout_3574+FA_out_3576+FA_cout_3589;
  assign {FA_cout_3716,FA_out_3716}=FA_cout_3576+FA_out_3578+FA_cout_3591;
  assign {FA_cout_3717,FA_out_3717}=FA_cout_3578+FA_out_3580+FA_cout_3593;
  assign {FA_cout_3718,FA_out_3718}=FA_cout_3580+FA_out_3582+HA_cout_223;
  assign {FA_cout_3719,FA_out_3719}=FA_cout_3582+FA_out_3584+HA_cout_224;
  assign {FA_cout_3720,FA_out_3720}=FA_cout_3584+FA_out_3586+HA_cout_225;
  assign {FA_cout_3721,FA_out_3721}=FA_cout_3586+FA_out_3588+HA_cout_226;
  assign {FA_cout_3722,FA_out_3722}=FA_cout_3588+FA_out_3590+FA_out_3415;
  assign {FA_cout_3723,FA_out_3723}=FA_cout_3590+FA_out_3592+FA_out_3419;
  assign {FA_cout_3724,FA_out_3724}=FA_cout_3592+FA_out_3594+FA_out_3423;
  assign {FA_cout_3725,FA_out_3725}=FA_cout_3594+FA_out_3595+FA_out_3427;
  assign {FA_cout_3726,FA_out_3726}=FA_cout_3595+FA_out_3596+FA_out_3431;
  assign {FA_cout_3727,FA_out_3727}=FA_cout_3596+FA_out_3597+FA_out_3435;
  assign {FA_cout_3728,FA_out_3728}=FA_cout_3597+FA_out_3598+HA_out_186;
  assign {FA_cout_3729,FA_out_3729}=FA_cout_3598+FA_out_3606+FA_out_3152;
  assign {FA_cout_3730,FA_out_3730}=FA_cout_3622+FA_out_3623+HA_out_219;
  assign {FA_cout_3731,FA_out_3731}=FA_cout_3623+FA_out_3624+HA_out_220;
  assign {FA_cout_3732,FA_out_3732}=FA_cout_3624+FA_out_3625+HA_out_221;
  assign {FA_cout_3733,FA_out_3733}=FA_cout_3625+FA_out_3626+HA_out_222;
  assign {FA_cout_3734,FA_out_3734}=FA_cout_3626+FA_out_3627+FA_out_3505;
  assign {FA_cout_3735,FA_out_3735}=FA_cout_3627+FA_out_3628+FA_out_3506;
  assign {FA_cout_3736,FA_out_3736}=FA_cout_3628+FA_out_3629+FA_out_3507;
  assign {FA_cout_3737,FA_out_3737}=FA_cout_3629+FA_out_3630+FA_out_3508;
  assign {FA_cout_3738,FA_out_3738}=FA_cout_3630+FA_out_3631+FA_out_3509;
  assign {FA_cout_3739,FA_out_3739}=FA_cout_3631+FA_out_3632+FA_out_3510;
  assign {FA_cout_3740,FA_out_3740}=FA_cout_3632+FA_out_3633+FA_out_3511;
  assign {FA_cout_3741,FA_out_3741}=FA_cout_3633+FA_out_3634+FA_out_3512;
  assign {FA_cout_3742,FA_out_3742}=FA_cout_3634+FA_out_3635+FA_out_3513;
  assign {FA_cout_3743,FA_out_3743}=FA_cout_3635+FA_out_3636+HA_out_277;
  assign {FA_cout_3744,FA_out_3744}=FA_cout_3636+FA_out_3637+HA_cout_277;
  assign {FA_cout_3745,FA_out_3745}=FA_cout_3637+FA_out_3638+HA_cout_278;
  assign {FA_cout_3746,FA_out_3746}=FA_cout_3638+FA_out_3639+HA_cout_279;
  assign {FA_cout_3747,FA_out_3747}=FA_cout_3639+FA_out_3640+HA_cout_280;
  assign {FA_cout_3748,FA_out_3748}=FA_cout_3640+FA_out_3641+HA_cout_281;
  assign {FA_cout_3749,FA_out_3749}=FA_cout_3641+FA_out_3642+HA_cout_282;
  assign {FA_cout_3750,FA_out_3750}=FA_cout_3642+FA_out_3643+HA_cout_283;
  assign {FA_cout_3751,FA_out_3751}=FA_cout_3643+FA_out_3644+HA_cout_284;
  assign {FA_cout_3752,FA_out_3752}=FA_cout_3644+FA_out_3645+FA_cout_3669;
  assign {FA_cout_3753,FA_out_3753}=FA_cout_3645+FA_out_3646+FA_cout_3670;
  assign {FA_cout_3754,FA_out_3754}=FA_cout_3646+FA_out_3647+FA_cout_3671;
  assign {FA_cout_3755,FA_out_3755}=FA_cout_3647+FA_out_3648+FA_cout_3672;
  assign {FA_cout_3756,FA_out_3756}=FA_cout_3648+FA_out_3649+FA_cout_3673;
  assign {FA_cout_3757,FA_out_3757}=FA_cout_3649+FA_out_3650+FA_cout_3674;
  assign {FA_cout_3758,FA_out_3758}=FA_cout_3650+FA_out_3651+FA_cout_3675;
  assign {FA_cout_3759,FA_out_3759}=FA_cout_3651+FA_out_3652+FA_cout_3676;
  assign {FA_cout_3760,FA_out_3760}=FA_cout_3652+FA_out_3653+FA_cout_3677;
  assign {FA_cout_3761,FA_out_3761}=FA_cout_3653+FA_out_3654+FA_cout_3678;
  assign {FA_cout_3762,FA_out_3762}=FA_cout_3654+FA_out_3655+FA_cout_3679;
  assign {FA_cout_3763,FA_out_3763}=FA_cout_3655+FA_out_3656+FA_cout_3680;
  assign {FA_cout_3764,FA_out_3764}=FA_cout_3656+FA_out_3657+FA_cout_3681;
  assign {FA_cout_3765,FA_out_3765}=FA_cout_3657+FA_out_3658+FA_cout_3682;
  assign {FA_cout_3766,FA_out_3766}=FA_cout_3658+FA_out_3659+FA_cout_3683;
  assign {FA_cout_3767,FA_out_3767}=FA_cout_3659+FA_out_3660+FA_cout_3684;
  assign {FA_cout_3768,FA_out_3768}=FA_cout_3660+FA_out_3661+FA_cout_3685;
  assign {FA_cout_3769,FA_out_3769}=FA_cout_3661+FA_out_3662+FA_cout_3687;
  assign {FA_cout_3770,FA_out_3770}=FA_cout_3662+FA_out_3663+FA_cout_3689;
  assign {FA_cout_3771,FA_out_3771}=FA_cout_3663+FA_out_3664+FA_cout_3691;
  assign {FA_cout_3772,FA_out_3772}=FA_cout_3664+FA_out_3665+FA_cout_3693;
  assign {FA_cout_3773,FA_out_3773}=FA_cout_3665+FA_out_3666+FA_cout_3695;
  assign {FA_cout_3774,FA_out_3774}=FA_cout_3666+FA_out_3667+FA_cout_3697;
  assign {FA_cout_3775,FA_out_3775}=FA_cout_3667+FA_out_3668+FA_cout_3699;
  assign {FA_cout_3776,FA_out_3776}=FA_cout_3668+FA_out_3686+FA_cout_3701;
  assign {FA_cout_3777,FA_out_3777}=FA_cout_3686+FA_out_3688+FA_cout_3703;
  assign {FA_cout_3778,FA_out_3778}=FA_cout_3688+FA_out_3690+FA_cout_3705;
  assign {FA_cout_3779,FA_out_3779}=FA_cout_3690+FA_out_3692+FA_cout_3707;
  assign {FA_cout_3780,FA_out_3780}=FA_cout_3692+FA_out_3694+FA_cout_3709;
  assign {FA_cout_3781,FA_out_3781}=FA_cout_3694+FA_out_3696+HA_cout_285;
  assign {FA_cout_3782,FA_out_3782}=FA_cout_3696+FA_out_3698+HA_cout_286;
  assign {FA_cout_3783,FA_out_3783}=FA_cout_3698+FA_out_3700+HA_cout_287;
  assign {FA_cout_3784,FA_out_3784}=FA_cout_3700+FA_out_3702+HA_cout_288;
  assign {FA_cout_3785,FA_out_3785}=FA_cout_3702+FA_out_3704+HA_cout_289;
  assign {FA_cout_3786,FA_out_3786}=FA_cout_3704+FA_out_3706+HA_cout_290;
  assign {FA_cout_3787,FA_out_3787}=FA_cout_3706+FA_out_3708+FA_out_3579;
  assign {FA_cout_3788,FA_out_3788}=FA_cout_3708+FA_out_3710+FA_out_3581;
  assign {FA_cout_3789,FA_out_3789}=FA_cout_3710+FA_out_3711+FA_out_3583;
  assign {FA_cout_3790,FA_out_3790}=FA_cout_3711+FA_out_3712+FA_out_3585;
  assign {FA_cout_3791,FA_out_3791}=FA_cout_3712+FA_out_3713+FA_out_3587;
  assign {FA_cout_3792,FA_out_3792}=FA_cout_3713+FA_out_3714+FA_out_3589;
  assign {FA_cout_3793,FA_out_3793}=FA_cout_3714+FA_out_3715+FA_out_3591;
  assign {FA_cout_3794,FA_out_3794}=FA_cout_3715+FA_out_3716+FA_out_3593;
  assign {FA_cout_3795,FA_out_3795}=FA_cout_3716+FA_out_3717+HA_out_223;
  assign {FA_cout_3796,FA_out_3796}=FA_cout_3717+FA_out_3718+HA_out_224;
  assign {FA_cout_3797,FA_out_3797}=FA_cout_3718+FA_out_3719+HA_out_225;
  assign {FA_cout_3798,FA_out_3798}=FA_cout_3719+FA_out_3720+HA_out_226;
  assign {FA_cout_3799,FA_out_3799}=FA_cout_3720+FA_out_3721+FA_out_3411;
  assign {FA_cout_3800,FA_out_3800}=REGS_1350+REGS_1413+REGS_1456;
  assign {FA_cout_3801,FA_out_3801}=REGS_1351+REGS_1414+REGS_1457;
  assign {FA_cout_3802,FA_out_3802}=REGS_1352+REGS_1415+REGS_1458;
  assign {FA_cout_3803,FA_out_3803}=REGS_1353+REGS_1416+REGS_1459;
  assign {FA_cout_3804,FA_out_3804}=REGS_1354+REGS_1417+REGS_1460;
  assign {FA_cout_3805,FA_out_3805}=REGS_1355+REGS_1418+REGS_1461;
  assign {FA_cout_3806,FA_out_3806}=REGS_1356+REGS_1419+REGS_1462;
  assign {FA_cout_3807,FA_out_3807}=REGS_1357+REGS_1420+REGS_1463;
  assign {FA_cout_3808,FA_out_3808}=REGS_1358+REGS_1421+REGS_1464;
  assign {FA_cout_3809,FA_out_3809}=REGS_1359+REGS_1422+REGS_1465;
  assign {FA_cout_3810,FA_out_3810}=REGS_1360+REGS_1423+REGS_1466;
  assign {FA_cout_3811,FA_out_3811}=REGS_1361+REGS_1424+REGS_1467;
  assign {FA_cout_3812,FA_out_3812}=REGS_1362+REGS_1425+REGS_1468;
  assign {FA_cout_3813,FA_out_3813}=REGS_1363+REGS_1426+REGS_1469;
  assign {FA_cout_3814,FA_out_3814}=REGS_1364+REGS_1427+REGS_1470;
  assign {FA_cout_3815,FA_out_3815}=REGS_1365+REGS_1428+REGS_1471;
  assign {FA_cout_3816,FA_out_3816}=REGS_1366+REGS_1429+REGS_1472;
  assign {FA_cout_3817,FA_out_3817}=REGS_1367+REGS_1430+REGS_1473;
  assign {FA_cout_3818,FA_out_3818}=REGS_1368+REGS_1431+REGS_1474;
  assign {FA_cout_3819,FA_out_3819}=REGS_1369+REGS_1432+REGS_1475;
  assign {FA_cout_3820,FA_out_3820}=REGS_1370+REGS_1433+REGS_1476;
  assign {FA_cout_3821,FA_out_3821}=REGS_1371+REGS_1434+REGS_1477;
  assign {FA_cout_3822,FA_out_3822}=REGS_1372+REGS_1435+REGS_1478;
  assign {FA_cout_3823,FA_out_3823}=REGS_1373+REGS_1436+REGS_1479;
  assign {FA_cout_3824,FA_out_3824}=REGS_1374+REGS_1437+REGS_1480;
  assign {FA_cout_3825,FA_out_3825}=REGS_1375+REGS_1438+REGS_1484;
  assign {FA_cout_3826,FA_out_3826}=REGS_1439+REGS_1440+REGS_1487;
  assign {FA_cout_3827,FA_out_3827}=REGS_1441+REGS_1442+REGS_1490;
  assign {FA_cout_3828,FA_out_3828}=REGS_1443+REGS_1444+REGS_1493;
  assign {FA_cout_3829,FA_out_3829}=REGS_1445+REGS_1446+REGS_1496;
  assign {FA_cout_3830,FA_out_3830}=REGS_1447+REGS_1448+REGS_1499;
  assign {FA_cout_3831,FA_out_3831}=REGS_1449+REGS_1450+REGS_1502;
  assign {FA_cout_3832,FA_out_3832}=REGS_1451+REGS_1452+REGS_1505;
  assign {FA_cout_3833,FA_out_3833}=REGS_1453+REGS_1454+REGS_1508;
  assign {FA_cout_3834,FA_out_3834}=REGS_1455+REGS_1481+REGS_1511;
  assign {FA_cout_3835,FA_out_3835}=REGS_1482+REGS_1485+REGS_1514;
  assign {FA_cout_3836,FA_out_3836}=REGS_1486+REGS_1488+REGS_1517;
  assign {FA_cout_3837,FA_out_3837}=REGS_1489+REGS_1491+REGS_1520;
  assign {FA_cout_3838,FA_out_3838}=REGS_1492+REGS_1494+REGS_1523;
  assign {FA_cout_3839,FA_out_3839}=REGS_1495+REGS_1497+REGS_1526;
  assign {FA_cout_3840,FA_out_3840}=REGS_1498+REGS_1500+REGS_1529;
  assign {FA_cout_3841,FA_out_3841}=REGS_1501+REGS_1503+REGS_1532;
  assign {FA_cout_3842,FA_out_3842}=REGS_1504+REGS_1506+REGS_1535;
  assign {FA_cout_3843,FA_out_3843}=FA_cout_3820+FA_out_3821+REGS_1483;
  assign {HA_cout_0,HA_out_0}=inp_0[1]+inp_1[0];
  assign {HA_cout_1,HA_out_1}=inp_3[1]+inp_4[0];
  assign {HA_cout_2,HA_out_2}=inp_6[1]+inp_7[0];
  assign {HA_cout_3,HA_out_3}=inp_9[1]+inp_10[0];
  assign {HA_cout_4,HA_out_4}=inp_12[1]+inp_13[0];
  assign {HA_cout_5,HA_out_5}=inp_15[1]+inp_16[0];
  assign {HA_cout_6,HA_out_6}=inp_18[1]+inp_19[0];
  assign {HA_cout_7,HA_out_7}=inp_21[1]+inp_22[0];
  assign {HA_cout_8,HA_out_8}=inp_24[1]+inp_25[0];
  assign {HA_cout_9,HA_out_9}=inp_27[1]+inp_28[0];
  assign {HA_cout_10,HA_out_10}=inp_30[1]+inp_31[0];
  assign {HA_cout_11,HA_out_11}=inp_33[1]+inp_34[0];
  assign {HA_cout_12,HA_out_12}=inp_36[1]+inp_37[0];
  assign {HA_cout_13,HA_out_13}=inp_39[1]+inp_40[0];
  assign {HA_cout_14,HA_out_14}=inp_42[1]+inp_43[0];
  assign {HA_cout_15,HA_out_15}=inp_45[1]+inp_46[0];
  assign {HA_cout_16,HA_out_16}=inp_48[1]+inp_49[0];
  assign {HA_cout_17,HA_out_17}=inp_51[1]+inp_52[0];
  assign {HA_cout_18,HA_out_18}=inp_54[1]+inp_55[0];
  assign {HA_cout_19,HA_out_19}=inp_57[1]+inp_58[0];
  assign {HA_cout_20,HA_out_20}=inp_60[1]+inp_61[0];
  assign {HA_cout_21,HA_out_21}=inp_62[3]+inp_63[2];
  assign {HA_cout_22,HA_out_22}=inp_62[6]+inp_63[5];
  assign {HA_cout_23,HA_out_23}=inp_62[9]+inp_63[8];
  assign {HA_cout_24,HA_out_24}=inp_62[12]+inp_63[11];
  assign {HA_cout_25,HA_out_25}=inp_62[15]+inp_63[14];
  assign {HA_cout_26,HA_out_26}=inp_62[18]+inp_63[17];
  assign {HA_cout_27,HA_out_27}=inp_62[21]+inp_63[20];
  assign {HA_cout_28,HA_out_28}=inp_62[24]+inp_63[23];
  assign {HA_cout_29,HA_out_29}=inp_62[27]+inp_63[26];
  assign {HA_cout_30,HA_out_30}=inp_62[30]+inp_63[29];
  assign {HA_cout_31,HA_out_31}=inp_62[33]+inp_63[32];
  assign {HA_cout_32,HA_out_32}=inp_62[36]+inp_63[35];
  assign {HA_cout_33,HA_out_33}=inp_62[39]+inp_63[38];
  assign {HA_cout_34,HA_out_34}=inp_62[42]+inp_63[41];
  assign {HA_cout_35,HA_out_35}=inp_62[45]+inp_63[44];
  assign {HA_cout_36,HA_out_36}=inp_62[48]+inp_63[47];
  assign {HA_cout_37,HA_out_37}=inp_62[51]+inp_63[50];
  assign {HA_cout_38,HA_out_38}=inp_62[54]+inp_63[53];
  assign {HA_cout_39,HA_out_39}=inp_62[57]+inp_63[56];
  assign {HA_cout_40,HA_out_40}=inp_62[60]+inp_63[59];
  assign {HA_cout_41,HA_out_41}=inp_62[63]+inp_63[62];
  assign {HA_cout_42,HA_out_42}=HA_cout_0+FA_out_0;
  assign {HA_cout_43,HA_out_43}=FA_out_65+inp_6[0];
  assign {HA_cout_44,HA_out_44}=FA_out_66+HA_out_2;
  assign {HA_cout_45,HA_out_45}=HA_cout_3+FA_out_192;
  assign {HA_cout_46,HA_out_46}=FA_out_257+inp_15[0];
  assign {HA_cout_47,HA_out_47}=FA_out_258+HA_out_5;
  assign {HA_cout_48,HA_out_48}=HA_cout_6+FA_out_384;
  assign {HA_cout_49,HA_out_49}=FA_out_449+inp_24[0];
  assign {HA_cout_50,HA_out_50}=FA_out_450+HA_out_8;
  assign {HA_cout_51,HA_out_51}=HA_cout_9+FA_out_576;
  assign {HA_cout_52,HA_out_52}=FA_out_641+inp_33[0];
  assign {HA_cout_53,HA_out_53}=FA_out_642+HA_out_11;
  assign {HA_cout_54,HA_out_54}=HA_cout_12+FA_out_768;
  assign {HA_cout_55,HA_out_55}=FA_out_833+inp_42[0];
  assign {HA_cout_56,HA_out_56}=FA_out_834+HA_out_14;
  assign {HA_cout_57,HA_out_57}=HA_cout_15+FA_out_960;
  assign {HA_cout_58,HA_out_58}=FA_out_1025+inp_51[0];
  assign {HA_cout_59,HA_out_59}=FA_out_1026+HA_out_17;
  assign {HA_cout_60,HA_out_60}=HA_cout_18+FA_out_1152;
  assign {HA_cout_61,HA_out_61}=FA_out_1217+inp_60[0];
  assign {HA_cout_62,HA_out_62}=FA_out_1218+HA_out_20;
  assign {HA_cout_63,HA_out_63}=FA_cout_1283+FA_out_1304;
  assign {HA_cout_64,HA_out_64}=FA_cout_1286+FA_out_1307;
  assign {HA_cout_65,HA_out_65}=FA_cout_1289+FA_out_1310;
  assign {HA_cout_66,HA_out_66}=FA_cout_1292+FA_out_1313;
  assign {HA_cout_67,HA_out_67}=FA_cout_1295+FA_out_1316;
  assign {HA_cout_68,HA_out_68}=FA_cout_1298+FA_out_1319;
  assign {HA_cout_69,HA_out_69}=FA_cout_1301+FA_out_1322;
  assign {HA_cout_70,HA_out_70}=FA_cout_1304+HA_out_23;
  assign {HA_cout_71,HA_out_71}=FA_cout_1307+HA_out_26;
  assign {HA_cout_72,HA_out_72}=FA_cout_1310+HA_out_29;
  assign {HA_cout_73,HA_out_73}=FA_cout_1313+HA_out_32;
  assign {HA_cout_74,HA_out_74}=FA_cout_1316+HA_out_35;
  assign {HA_cout_75,HA_out_75}=FA_cout_1319+HA_out_38;
  assign {HA_cout_76,HA_out_76}=FA_cout_1322+HA_out_41;
  assign {HA_cout_77,HA_out_77}=HA_cout_23+inp_63[9];
  assign {HA_cout_78,HA_out_78}=HA_cout_26+inp_63[18];
  assign {HA_cout_79,HA_out_79}=HA_cout_29+inp_63[27];
  assign {HA_cout_80,HA_out_80}=HA_cout_32+inp_63[36];
  assign {HA_cout_81,HA_out_81}=HA_cout_35+inp_63[45];
  assign {HA_cout_82,HA_out_82}=HA_cout_38+inp_63[54];
  assign {HA_cout_83,HA_out_83}=HA_cout_41+inp_63[63];
  assign {HA_cout_84,HA_out_84}=HA_cout_42+FA_out_1323;
  assign {HA_cout_85,HA_out_85}=FA_cout_1323+FA_out_1324;
  assign {HA_cout_86,HA_out_86}=FA_out_1389+inp_9[0];
  assign {HA_cout_87,HA_out_87}=FA_out_1390+HA_out_3;
  assign {HA_cout_88,HA_out_88}=FA_out_1391+HA_out_45;
  assign {HA_cout_89,HA_out_89}=HA_cout_46+HA_out_47;
  assign {HA_cout_90,HA_out_90}=HA_cout_47+FA_out_1518;
  assign {HA_cout_91,HA_out_91}=FA_out_1587+FA_out_448;
  assign {HA_cout_92,HA_out_92}=FA_out_1588+HA_out_49;
  assign {HA_cout_93,HA_out_93}=HA_cout_51+FA_out_1716;
  assign {HA_cout_94,HA_out_94}=FA_cout_1716+FA_out_1717;
  assign {HA_cout_95,HA_out_95}=FA_out_1779+inp_36[0];
  assign {HA_cout_96,HA_out_96}=FA_out_1780+HA_out_12;
  assign {HA_cout_97,HA_out_97}=FA_out_1781+HA_out_54;
  assign {HA_cout_98,HA_out_98}=HA_cout_55+HA_out_56;
  assign {HA_cout_99,HA_out_99}=HA_cout_56+FA_out_1908;
  assign {HA_cout_100,HA_out_100}=FA_out_1980+FA_out_1024;
  assign {HA_cout_101,HA_out_101}=FA_out_1981+HA_out_58;
  assign {HA_cout_102,HA_out_102}=HA_cout_60+FA_out_2109;
  assign {HA_cout_103,HA_out_103}=FA_cout_2109+FA_out_2110;
  assign {HA_cout_104,HA_out_104}=FA_out_2173+HA_out_25;
  assign {HA_cout_105,HA_out_105}=FA_cout_2174+FA_out_2188;
  assign {HA_cout_106,HA_out_106}=FA_out_2176+HA_cout_79;
  assign {HA_cout_107,HA_out_107}=FA_out_2179+HA_out_34;
  assign {HA_cout_108,HA_out_108}=FA_cout_2180+FA_out_2194;
  assign {HA_cout_109,HA_out_109}=FA_out_2182+HA_cout_82;
  assign {HA_cout_110,HA_out_110}=FA_out_2169+inp_63[0];
  assign {HA_cout_111,HA_out_111}=FA_cout_2185+HA_out_63;
  assign {HA_cout_112,HA_out_112}=FA_out_2187+inp_63[15];
  assign {HA_cout_113,HA_out_113}=FA_cout_2188+FA_out_2200;
  assign {HA_cout_114,HA_out_114}=FA_cout_2191+HA_out_66;
  assign {HA_cout_115,HA_out_115}=FA_out_2193+inp_63[42];
  assign {HA_cout_116,HA_out_116}=FA_cout_2194+FA_out_2203;
  assign {HA_cout_117,HA_out_117}=FA_cout_2197+HA_out_69;
  assign {HA_cout_118,HA_out_118}=HA_cout_63+HA_out_70;
  assign {HA_cout_119,HA_out_119}=FA_cout_2200+FA_out_1309;
  assign {HA_cout_120,HA_out_120}=HA_cout_66+HA_out_73;
  assign {HA_cout_121,HA_out_121}=FA_cout_2203+FA_out_1318;
  assign {HA_cout_122,HA_out_122}=HA_cout_69+HA_out_76;
  assign {HA_cout_123,HA_out_123}=HA_cout_70+HA_out_77;
  assign {HA_cout_124,HA_out_124}=HA_cout_73+HA_out_80;
  assign {HA_cout_125,HA_out_125}=HA_cout_76+HA_out_83;
  assign {HA_cout_126,HA_out_126}=REGS_4+REGS_67;
  assign {HA_cout_127,HA_out_127}=REGS_5+REGS_68;
  assign {HA_cout_128,HA_out_128}=REGS_6+REGS_69;
  assign {HA_cout_129,HA_out_129}=REGS_203+REGS_283;
  assign {HA_cout_130,HA_out_130}=REGS_204+REGS_284;
  assign {HA_cout_131,HA_out_131}=REGS_205+REGS_285;
  assign {HA_cout_132,HA_out_132}=REGS_422+REGS_471;
  assign {HA_cout_133,HA_out_133}=REGS_423+REGS_472;
  assign {HA_cout_134,HA_out_134}=REGS_424+REGS_473;
  assign {HA_cout_135,HA_out_135}=REGS_620+REGS_692;
  assign {HA_cout_136,HA_out_136}=REGS_621+REGS_693;
  assign {HA_cout_137,HA_out_137}=REGS_622+REGS_694;
  assign {HA_cout_138,HA_out_138}=REGS_851+REGS_886;
  assign {HA_cout_139,HA_out_139}=REGS_852+REGS_887;
  assign {HA_cout_140,HA_out_140}=REGS_853+REGS_888;
  assign {HA_cout_141,HA_out_141}=REGS_854+REGS_889;
  assign {HA_cout_142,HA_out_142}=REGS_1014+REGS_1138;
  assign {HA_cout_143,HA_out_143}=REGS_1015+REGS_1139;
  assign {HA_cout_144,HA_out_144}=REGS_1016+REGS_1140;
  assign {HA_cout_145,HA_out_145}=REGS_1017+REGS_1141;
  assign {HA_cout_146,HA_out_146}=REGS_1160+REGS_1185;
  assign {HA_cout_147,HA_out_147}=REGS_1163+REGS_1303;
  assign {HA_cout_148,HA_out_148}=REGS_1183+REGS_1275;
  assign {HA_cout_149,HA_out_149}=REGS_1186+REGS_1203;
  assign {HA_cout_150,HA_out_150}=REGS_1198+REGS_1215;
  assign {HA_cout_151,HA_out_151}=REGS_1201+REGS_1288;
  assign {HA_cout_152,HA_out_152}=REGS_1204+REGS_1221;
  assign {HA_cout_153,HA_out_153}=REGS_1210+REGS_1227;
  assign {HA_cout_154,HA_out_154}=REGS_1216+REGS_1233;
  assign {HA_cout_155,HA_out_155}=REGS_1222+REGS_1239;
  assign {HA_cout_156,HA_out_156}=REGS_1228+REGS_1245;
  assign {HA_cout_157,HA_out_157}=REGS_1234+REGS_1256;
  assign {HA_cout_158,HA_out_158}=REGS_1240+REGS_1261;
  assign {HA_cout_159,HA_out_159}=REGS_1246+REGS_1266;
  assign {HA_cout_160,HA_out_160}=REGS_1250+REGS_1268;
  assign {HA_cout_161,HA_out_161}=REGS_1257+REGS_1273;
  assign {HA_cout_162,HA_out_162}=REGS_1262+REGS_1278;
  assign {HA_cout_163,HA_out_163}=REGS_1267+REGS_1282;
  assign {HA_cout_164,HA_out_164}=REGS_1274+REGS_1297;
  assign {HA_cout_165,HA_out_165}=REGS_1283+REGS_1293;
  assign {HA_cout_166,HA_out_166}=REGS_1294+REGS_1301;
  assign {HA_cout_167,HA_out_167}=HA_cout_126+HA_out_127;
  assign {HA_cout_168,HA_out_168}=HA_cout_127+HA_out_128;
  assign {HA_cout_169,HA_out_169}=HA_cout_128+FA_out_2792;
  assign {HA_cout_170,HA_out_170}=FA_cout_2792+FA_out_2793;
  assign {HA_cout_171,HA_out_171}=FA_cout_2793+FA_out_2794;
  assign {HA_cout_172,HA_out_172}=FA_out_2861+REGS_419;
  assign {HA_cout_173,HA_out_173}=FA_out_2862+REGS_420;
  assign {HA_cout_174,HA_out_174}=FA_out_2863+REGS_421;
  assign {HA_cout_175,HA_out_175}=FA_out_2864+HA_out_132;
  assign {HA_cout_176,HA_out_176}=HA_cout_135+HA_out_136;
  assign {HA_cout_177,HA_out_177}=HA_cout_136+HA_out_137;
  assign {HA_cout_178,HA_out_178}=HA_cout_137+FA_out_2998;
  assign {HA_cout_179,HA_out_179}=FA_cout_2998+FA_out_2999;
  assign {HA_cout_180,HA_out_180}=FA_cout_2999+FA_out_3000;
  assign {HA_cout_181,HA_out_181}=FA_cout_3000+FA_out_3001;
  assign {HA_cout_182,HA_out_182}=FA_out_3078+REGS_1011;
  assign {HA_cout_183,HA_out_183}=FA_out_3079+REGS_1012;
  assign {HA_cout_184,HA_out_184}=FA_out_3080+REGS_1013;
  assign {HA_cout_185,HA_out_185}=FA_out_3081+HA_out_142;
  assign {HA_cout_186,HA_out_186}=FA_out_3146+REGS_1299;
  assign {HA_cout_187,HA_out_187}=FA_out_3149+REGS_1195;
  assign {HA_cout_188,HA_out_188}=FA_cout_3150+FA_out_3156;
  assign {HA_cout_189,HA_out_189}=FA_out_3155+REGS_1213;
  assign {HA_cout_190,HA_out_190}=FA_cout_3156+FA_out_3162;
  assign {HA_cout_191,HA_out_191}=FA_out_3161+REGS_1231;
  assign {HA_cout_192,HA_out_192}=FA_cout_3162+FA_out_3168;
  assign {HA_cout_193,HA_out_193}=FA_out_3167+REGS_1254;
  assign {HA_cout_194,HA_out_194}=FA_cout_3168+FA_out_3174;
  assign {HA_cout_195,HA_out_195}=FA_out_3173+REGS_1272;
  assign {HA_cout_196,HA_out_196}=FA_cout_3174+FA_out_3180;
  assign {HA_cout_197,HA_out_197}=FA_cout_3177+FA_out_3181;
  assign {HA_cout_198,HA_out_198}=FA_cout_3180+HA_out_148;
  assign {HA_cout_199,HA_out_199}=FA_cout_3181+FA_out_3183;
  assign {HA_cout_200,HA_out_200}=HA_cout_148+HA_out_151;
  assign {HA_cout_201,HA_out_201}=FA_cout_3183+HA_out_153;
  assign {HA_cout_202,HA_out_202}=HA_cout_151+REGS_1219;
  assign {HA_cout_203,HA_out_203}=HA_cout_153+HA_out_156;
  assign {HA_cout_204,HA_out_204}=HA_cout_156+HA_out_159;
  assign {HA_cout_205,HA_out_205}=HA_cout_159+HA_out_163;
  assign {HA_cout_206,HA_out_206}=HA_cout_160+REGS_1251;
  assign {HA_cout_207,HA_out_207}=HA_cout_163+HA_out_165;
  assign {HA_cout_208,HA_out_208}=HA_cout_165+HA_out_166;
  assign {HA_cout_209,HA_out_209}=HA_cout_167+HA_out_168;
  assign {HA_cout_210,HA_out_210}=HA_cout_168+HA_out_169;
  assign {HA_cout_211,HA_out_211}=HA_cout_169+HA_out_170;
  assign {HA_cout_212,HA_out_212}=HA_cout_170+HA_out_171;
  assign {HA_cout_213,HA_out_213}=HA_cout_171+FA_out_3184;
  assign {HA_cout_214,HA_out_214}=FA_cout_3184+FA_out_3185;
  assign {HA_cout_215,HA_out_215}=FA_cout_3185+FA_out_3186;
  assign {HA_cout_216,HA_out_216}=FA_cout_3186+FA_out_3187;
  assign {HA_cout_217,HA_out_217}=FA_cout_3187+FA_out_3188;
  assign {HA_cout_218,HA_out_218}=FA_out_3254+REGS_617;
  assign {HA_cout_219,HA_out_219}=FA_out_3255+REGS_618;
  assign {HA_cout_220,HA_out_220}=FA_out_3256+REGS_619;
  assign {HA_cout_221,HA_out_221}=FA_out_3257+HA_out_135;
  assign {HA_cout_222,HA_out_222}=FA_out_3258+HA_out_176;
  assign {HA_cout_223,HA_out_223}=FA_out_3386+REGS_1259;
  assign {HA_cout_224,HA_out_224}=FA_out_3389+REGS_1276;
  assign {HA_cout_225,HA_out_225}=FA_out_3392+REGS_1289;
  assign {HA_cout_226,HA_out_226}=FA_out_3395+REGS_1298;
  assign {HA_cout_227,HA_out_227}=HA_cout_182+HA_out_183;
  assign {HA_cout_228,HA_out_228}=HA_cout_183+HA_out_184;
  assign {HA_cout_229,HA_out_229}=HA_cout_184+HA_out_185;
  assign {HA_cout_230,HA_out_230}=HA_cout_185+FA_out_3397;
  assign {HA_cout_231,HA_out_231}=FA_cout_3397+FA_out_3398;
  assign {HA_cout_232,HA_out_232}=FA_cout_3398+FA_out_3399;
  assign {HA_cout_233,HA_out_233}=FA_cout_3399+FA_out_3400;
  assign {HA_cout_234,HA_out_234}=FA_cout_3400+FA_out_3401;
  assign {HA_cout_235,HA_out_235}=FA_cout_3401+FA_out_3402;
  assign {HA_cout_236,HA_out_236}=FA_cout_3409+FA_out_3413;
  assign {HA_cout_237,HA_out_237}=FA_cout_3413+FA_out_3417;
  assign {HA_cout_238,HA_out_238}=FA_cout_3417+FA_out_3421;
  assign {HA_cout_239,HA_out_239}=FA_cout_3421+FA_out_3425;
  assign {HA_cout_240,HA_out_240}=FA_cout_3425+FA_out_3429;
  assign {HA_cout_241,HA_out_241}=FA_cout_3429+FA_out_3433;
  assign {HA_cout_242,HA_out_242}=FA_cout_3433+FA_out_3437;
  assign {HA_cout_243,HA_out_243}=FA_cout_3437+HA_out_187;
  assign {HA_cout_244,HA_out_244}=FA_cout_3439+FA_out_3440;
  assign {HA_cout_245,HA_out_245}=HA_cout_187+HA_out_189;
  assign {HA_cout_246,HA_out_246}=FA_cout_3440+FA_out_3441;
  assign {HA_cout_247,HA_out_247}=HA_cout_189+HA_out_191;
  assign {HA_cout_248,HA_out_248}=FA_cout_3441+FA_out_3442;
  assign {HA_cout_249,HA_out_249}=HA_cout_191+HA_out_193;
  assign {HA_cout_250,HA_out_250}=FA_cout_3442+FA_out_3443;
  assign {HA_cout_251,HA_out_251}=HA_cout_193+HA_out_195;
  assign {HA_cout_252,HA_out_252}=FA_cout_3443+HA_out_197;
  assign {HA_cout_253,HA_out_253}=HA_cout_195+FA_out_3179;
  assign {HA_cout_254,HA_out_254}=HA_cout_197+HA_out_199;
  assign {HA_cout_255,HA_out_255}=HA_cout_199+HA_out_201;
  assign {HA_cout_256,HA_out_256}=HA_cout_201+HA_out_203;
  assign {HA_cout_257,HA_out_257}=HA_cout_203+HA_out_204;
  assign {HA_cout_258,HA_out_258}=HA_cout_204+HA_out_205;
  assign {HA_cout_259,HA_out_259}=HA_cout_205+HA_out_207;
  assign {HA_cout_260,HA_out_260}=HA_cout_207+HA_out_208;
  assign {HA_cout_261,HA_out_261}=HA_cout_208+HA_cout_166;
  assign {HA_cout_262,HA_out_262}=HA_cout_209+HA_out_210;
  assign {HA_cout_263,HA_out_263}=HA_cout_210+HA_out_211;
  assign {HA_cout_264,HA_out_264}=HA_cout_211+HA_out_212;
  assign {HA_cout_265,HA_out_265}=HA_cout_212+HA_out_213;
  assign {HA_cout_266,HA_out_266}=HA_cout_213+HA_out_214;
  assign {HA_cout_267,HA_out_267}=HA_cout_214+HA_out_215;
  assign {HA_cout_268,HA_out_268}=HA_cout_215+HA_out_216;
  assign {HA_cout_269,HA_out_269}=HA_cout_216+HA_out_217;
  assign {HA_cout_270,HA_out_270}=HA_cout_217+FA_out_3444;
  assign {HA_cout_271,HA_out_271}=FA_cout_3444+FA_out_3445;
  assign {HA_cout_272,HA_out_272}=FA_cout_3445+FA_out_3446;
  assign {HA_cout_273,HA_out_273}=FA_cout_3446+FA_out_3447;
  assign {HA_cout_274,HA_out_274}=FA_cout_3447+FA_out_3448;
  assign {HA_cout_275,HA_out_275}=FA_cout_3448+FA_out_3449;
  assign {HA_cout_276,HA_out_276}=FA_cout_3449+FA_out_3450;
  assign {HA_cout_277,HA_out_277}=FA_out_3514+HA_out_139;
  assign {HA_cout_278,HA_out_278}=FA_out_3515+HA_out_140;
  assign {HA_cout_279,HA_out_279}=FA_out_3516+HA_out_141;
  assign {HA_cout_280,HA_out_280}=FA_out_3517+FA_out_3075;
  assign {HA_cout_281,HA_out_281}=FA_out_3518+FA_out_3076;
  assign {HA_cout_282,HA_out_282}=FA_out_3519+FA_out_3077;
  assign {HA_cout_283,HA_out_283}=FA_out_3520+HA_out_182;
  assign {HA_cout_284,HA_out_284}=FA_out_3521+HA_out_227;
  assign {HA_cout_285,HA_out_285}=FA_out_3565+HA_out_150;
  assign {HA_cout_286,HA_out_286}=FA_out_3567+HA_out_154;
  assign {HA_cout_287,HA_out_287}=FA_out_3569+HA_out_157;
  assign {HA_cout_288,HA_out_288}=FA_out_3571+HA_out_161;
  assign {HA_cout_289,HA_out_289}=FA_out_3573+HA_out_164;
  assign {HA_cout_290,HA_out_290}=FA_out_3575+REGS_1302;
  assign {HA_cout_291,HA_out_291}=FA_cout_3606+FA_out_3607;
  assign {HA_cout_292,HA_out_292}=FA_cout_3607+FA_out_3608;
  assign {HA_cout_293,HA_out_293}=FA_cout_3608+FA_out_3609;
  assign {HA_cout_294,HA_out_294}=FA_cout_3609+FA_out_3610;
  assign {HA_cout_295,HA_out_295}=FA_cout_3610+FA_out_3611;
  assign {HA_cout_296,HA_out_296}=FA_cout_3611+FA_out_3612;
  assign {HA_cout_297,HA_out_297}=FA_cout_3612+HA_out_244;
  assign {HA_cout_298,HA_out_298}=HA_cout_244+HA_out_246;
  assign {HA_cout_299,HA_out_299}=HA_cout_246+HA_out_248;
  assign {HA_cout_300,HA_out_300}=HA_cout_248+HA_out_250;
  assign {HA_cout_301,HA_out_301}=HA_cout_250+HA_out_252;
  assign {HA_cout_302,HA_out_302}=HA_cout_252+HA_out_254;
  assign {HA_cout_303,HA_out_303}=HA_cout_254+HA_out_255;
  assign {HA_cout_304,HA_out_304}=HA_cout_255+HA_out_256;
  assign {HA_cout_305,HA_out_305}=HA_cout_256+HA_out_257;
  assign {HA_cout_306,HA_out_306}=HA_cout_257+HA_out_258;
  assign {HA_cout_307,HA_out_307}=HA_cout_258+HA_out_259;
  assign {HA_cout_308,HA_out_308}=HA_cout_259+HA_out_260;
  assign {HA_cout_309,HA_out_309}=HA_cout_260+HA_out_261;
  assign {HA_cout_310,HA_out_310}=HA_cout_262+HA_out_263;
  assign {HA_cout_311,HA_out_311}=HA_cout_263+HA_out_264;
  assign {HA_cout_312,HA_out_312}=HA_cout_264+HA_out_265;
  assign {HA_cout_313,HA_out_313}=HA_cout_265+HA_out_266;
  assign {HA_cout_314,HA_out_314}=HA_cout_266+HA_out_267;
  assign {HA_cout_315,HA_out_315}=HA_cout_267+HA_out_268;
  assign {HA_cout_316,HA_out_316}=HA_cout_268+HA_out_269;
  assign {HA_cout_317,HA_out_317}=HA_cout_269+HA_out_270;
  assign {HA_cout_318,HA_out_318}=HA_cout_270+HA_out_271;
  assign {HA_cout_319,HA_out_319}=HA_cout_271+HA_out_272;
  assign {HA_cout_320,HA_out_320}=HA_cout_272+HA_out_273;
  assign {HA_cout_321,HA_out_321}=HA_cout_273+HA_out_274;
  assign {HA_cout_322,HA_out_322}=HA_cout_274+HA_out_275;
  assign {HA_cout_323,HA_out_323}=HA_cout_275+HA_out_276;
  assign {HA_cout_324,HA_out_324}=HA_cout_276+FA_out_3613;
  assign {HA_cout_325,HA_out_325}=FA_cout_3613+FA_out_3614;
  assign {HA_cout_326,HA_out_326}=FA_cout_3614+FA_out_3615;
  assign {HA_cout_327,HA_out_327}=FA_cout_3615+FA_out_3616;
  assign {HA_cout_328,HA_out_328}=FA_cout_3616+FA_out_3617;
  assign {HA_cout_329,HA_out_329}=FA_cout_3617+FA_out_3618;
  assign {HA_cout_330,HA_out_330}=FA_cout_3618+FA_out_3619;
  assign {HA_cout_331,HA_out_331}=FA_cout_3619+FA_out_3620;
  assign {HA_cout_332,HA_out_332}=FA_cout_3620+FA_out_3621;
  assign {HA_cout_333,HA_out_333}=FA_cout_3621+FA_out_3622;
  assign {HA_cout_334,HA_out_334}=FA_out_3682+REGS_1269;
  assign {HA_cout_335,HA_out_335}=FA_cout_3721+FA_out_3722;
  assign {HA_cout_336,HA_out_336}=FA_cout_3722+FA_out_3723;
  assign {HA_cout_337,HA_out_337}=FA_cout_3723+FA_out_3724;
  assign {HA_cout_338,HA_out_338}=FA_cout_3724+FA_out_3725;
  assign {HA_cout_339,HA_out_339}=FA_cout_3725+FA_out_3726;
  assign {HA_cout_340,HA_out_340}=FA_cout_3726+FA_out_3727;
  assign {HA_cout_341,HA_out_341}=FA_cout_3727+FA_out_3728;
  assign {HA_cout_342,HA_out_342}=FA_cout_3728+FA_out_3729;
  assign {HA_cout_343,HA_out_343}=FA_cout_3729+HA_out_291;
  assign {HA_cout_344,HA_out_344}=HA_cout_291+HA_out_292;
  assign {HA_cout_345,HA_out_345}=HA_cout_292+HA_out_293;
  assign {HA_cout_346,HA_out_346}=HA_cout_293+HA_out_294;
  assign {HA_cout_347,HA_out_347}=HA_cout_294+HA_out_295;
  assign {HA_cout_348,HA_out_348}=HA_cout_295+HA_out_296;
  assign {HA_cout_349,HA_out_349}=HA_cout_296+HA_out_297;
  assign {HA_cout_350,HA_out_350}=HA_cout_297+HA_out_298;
  assign {HA_cout_351,HA_out_351}=HA_cout_298+HA_out_299;
  assign {HA_cout_352,HA_out_352}=HA_cout_299+HA_out_300;
  assign {HA_cout_353,HA_out_353}=HA_cout_300+HA_out_301;
  assign {HA_cout_354,HA_out_354}=HA_cout_301+HA_out_302;
  assign {HA_cout_355,HA_out_355}=HA_cout_302+HA_out_303;
  assign {HA_cout_356,HA_out_356}=HA_cout_303+HA_out_304;
  assign {HA_cout_357,HA_out_357}=HA_cout_304+HA_out_305;
  assign {HA_cout_358,HA_out_358}=HA_cout_305+HA_out_306;
  assign {HA_cout_359,HA_out_359}=HA_cout_306+HA_out_307;
  assign {HA_cout_360,HA_out_360}=HA_cout_307+HA_out_308;
  assign {HA_cout_361,HA_out_361}=HA_cout_308+HA_out_309;
  assign {HA_cout_362,HA_out_362}=HA_cout_309+HA_cout_261;
  assign {HA_cout_363,HA_out_363}=REGS_1313+REGS_1376;
  assign {HA_cout_364,HA_out_364}=REGS_1314+REGS_1377;
  assign {HA_cout_365,HA_out_365}=REGS_1315+REGS_1378;
  assign {HA_cout_366,HA_out_366}=REGS_1316+REGS_1379;
  assign {HA_cout_367,HA_out_367}=REGS_1317+REGS_1380;
  assign {HA_cout_368,HA_out_368}=REGS_1318+REGS_1381;
  assign {HA_cout_369,HA_out_369}=REGS_1319+REGS_1382;
  assign {HA_cout_370,HA_out_370}=REGS_1320+REGS_1383;
  assign {HA_cout_371,HA_out_371}=REGS_1321+REGS_1384;
  assign {HA_cout_372,HA_out_372}=REGS_1322+REGS_1385;
  assign {HA_cout_373,HA_out_373}=REGS_1323+REGS_1386;
  assign {HA_cout_374,HA_out_374}=REGS_1324+REGS_1387;
  assign {HA_cout_375,HA_out_375}=REGS_1325+REGS_1388;
  assign {HA_cout_376,HA_out_376}=REGS_1326+REGS_1389;
  assign {HA_cout_377,HA_out_377}=REGS_1327+REGS_1390;
  assign {HA_cout_378,HA_out_378}=REGS_1328+REGS_1391;
  assign {HA_cout_379,HA_out_379}=REGS_1329+REGS_1392;
  assign {HA_cout_380,HA_out_380}=REGS_1330+REGS_1393;
  assign {HA_cout_381,HA_out_381}=REGS_1331+REGS_1394;
  assign {HA_cout_382,HA_out_382}=REGS_1332+REGS_1395;
  assign {HA_cout_383,HA_out_383}=REGS_1333+REGS_1396;
  assign {HA_cout_384,HA_out_384}=REGS_1334+REGS_1397;
  assign {HA_cout_385,HA_out_385}=REGS_1335+REGS_1398;
  assign {HA_cout_386,HA_out_386}=REGS_1336+REGS_1399;
  assign {HA_cout_387,HA_out_387}=REGS_1337+REGS_1400;
  assign {HA_cout_388,HA_out_388}=REGS_1338+REGS_1401;
  assign {HA_cout_389,HA_out_389}=REGS_1339+REGS_1402;
  assign {HA_cout_390,HA_out_390}=REGS_1340+REGS_1403;
  assign {HA_cout_391,HA_out_391}=REGS_1341+REGS_1404;
  assign {HA_cout_392,HA_out_392}=REGS_1342+REGS_1405;
  assign {HA_cout_393,HA_out_393}=REGS_1343+REGS_1406;
  assign {HA_cout_394,HA_out_394}=REGS_1344+REGS_1407;
  assign {HA_cout_395,HA_out_395}=REGS_1345+REGS_1408;
  assign {HA_cout_396,HA_out_396}=REGS_1346+REGS_1409;
  assign {HA_cout_397,HA_out_397}=REGS_1347+REGS_1410;
  assign {HA_cout_398,HA_out_398}=REGS_1348+REGS_1411;
  assign {HA_cout_399,HA_out_399}=REGS_1349+REGS_1412;
  assign {HA_cout_400,HA_out_400}=REGS_1507+REGS_1509;
  assign {HA_cout_401,HA_out_401}=REGS_1510+REGS_1512;
  assign {HA_cout_402,HA_out_402}=REGS_1513+REGS_1515;
  assign {HA_cout_403,HA_out_403}=REGS_1516+REGS_1518;
  assign {HA_cout_404,HA_out_404}=REGS_1519+REGS_1521;
  assign {HA_cout_405,HA_out_405}=REGS_1522+REGS_1524;
  assign {HA_cout_406,HA_out_406}=REGS_1525+REGS_1527;
  assign {HA_cout_407,HA_out_407}=REGS_1528+REGS_1530;
  assign {HA_cout_408,HA_out_408}=REGS_1531+REGS_1533;
  assign {HA_cout_409,HA_out_409}=REGS_1534+REGS_1536;
  assign {HA_cout_410,HA_out_410}=REGS_1537+REGS_1538;
  assign {HA_cout_411,HA_out_411}=REGS_1539+REGS_1540;
  assign {HA_cout_412,HA_out_412}=REGS_1541+REGS_1542;
  assign {HA_cout_413,HA_out_413}=REGS_1543+REGS_1544;
  assign {HA_cout_414,HA_out_414}=REGS_1545+REGS_1546;
  assign {HA_cout_415,HA_out_415}=REGS_1547+REGS_1548;
  assign {HA_cout_416,HA_out_416}=REGS_1549+REGS_1550;
  assign {HA_cout_417,HA_out_417}=REGS_1551+REGS_1552;
  assign {HA_cout_418,HA_out_418}=REGS_1553+REGS_1554;
  assign {HA_cout_419,HA_out_419}=REGS_1555+REGS_1556;
  assign {HA_cout_420,HA_out_420}=REGS_1557+REGS_1558;
  assign {HA_cout_421,HA_out_421}=REGS_1559+REGS_1560;
  assign {HA_cout_422,HA_out_422}=REGS_1561+REGS_1562;
  assign {HA_cout_423,HA_out_423}=REGS_1563+REGS_1564;
  assign {HA_cout_424,HA_out_424}=REGS_1565+REGS_1566;
  assign {HA_cout_425,HA_out_425}=REGS_1567+REGS_1568;
  assign {HA_cout_426,HA_out_426}=REGS_1569+REGS_1570;
  assign {HA_cout_427,HA_out_427}=REGS_1571+REGS_1572;
  assign {HA_cout_428,HA_out_428}=REGS_1573+REGS_1574;
  assign {HA_cout_429,HA_out_429}=REGS_1575+REGS_1576;
  assign {HA_cout_430,HA_out_430}=REGS_1577+REGS_1578;
  assign {HA_cout_431,HA_out_431}=REGS_1579+REGS_1580;
  assign {HA_cout_432,HA_out_432}=REGS_1581+REGS_1582;
  assign {HA_cout_433,HA_out_433}=REGS_1583+REGS_1584;
  assign {HA_cout_434,HA_out_434}=REGS_1585+REGS_1586;
  assign {HA_cout_435,HA_out_435}=REGS_1587+REGS_1588;
  assign {HA_cout_436,HA_out_436}=REGS_1589+REGS_1590;
  assign {HA_cout_437,HA_out_437}=REGS_1591+REGS_1592;
  assign {HA_cout_438,HA_out_438}=REGS_1593+REGS_1594;
  assign {HA_cout_439,HA_out_439}=REGS_1595+REGS_1596;
  assign {HA_cout_440,HA_out_440}=REGS_1597+REGS_1598;
  assign {HA_cout_441,HA_out_441}=HA_cout_363+HA_out_364;
  assign {HA_cout_442,HA_out_442}=HA_cout_364+HA_out_365;
  assign {HA_cout_443,HA_out_443}=HA_cout_365+HA_out_366;
  assign {HA_cout_444,HA_out_444}=HA_cout_366+HA_out_367;
  assign {HA_cout_445,HA_out_445}=HA_cout_367+HA_out_368;
  assign {HA_cout_446,HA_out_446}=HA_cout_368+HA_out_369;
  assign {HA_cout_447,HA_out_447}=HA_cout_369+HA_out_370;
  assign {HA_cout_448,HA_out_448}=HA_cout_370+HA_out_371;
  assign {HA_cout_449,HA_out_449}=HA_cout_371+HA_out_372;
  assign {HA_cout_450,HA_out_450}=HA_cout_372+HA_out_373;
  assign {HA_cout_451,HA_out_451}=HA_cout_373+HA_out_374;
  assign {HA_cout_452,HA_out_452}=HA_cout_374+HA_out_375;
  assign {HA_cout_453,HA_out_453}=HA_cout_375+HA_out_376;
  assign {HA_cout_454,HA_out_454}=HA_cout_376+HA_out_377;
  assign {HA_cout_455,HA_out_455}=HA_cout_377+HA_out_378;
  assign {HA_cout_456,HA_out_456}=HA_cout_378+HA_out_379;
  assign {HA_cout_457,HA_out_457}=HA_cout_379+HA_out_380;
  assign {HA_cout_458,HA_out_458}=HA_cout_380+HA_out_381;
  assign {HA_cout_459,HA_out_459}=HA_cout_381+HA_out_382;
  assign {HA_cout_460,HA_out_460}=HA_cout_382+HA_out_383;
  assign {HA_cout_461,HA_out_461}=HA_cout_383+HA_out_384;
  assign {HA_cout_462,HA_out_462}=HA_cout_384+HA_out_385;
  assign {HA_cout_463,HA_out_463}=HA_cout_385+HA_out_386;
  assign {HA_cout_464,HA_out_464}=HA_cout_386+HA_out_387;
  assign {HA_cout_465,HA_out_465}=HA_cout_387+HA_out_388;
  assign {HA_cout_466,HA_out_466}=HA_cout_388+HA_out_389;
  assign {HA_cout_467,HA_out_467}=HA_cout_389+HA_out_390;
  assign {HA_cout_468,HA_out_468}=HA_cout_390+HA_out_391;
  assign {HA_cout_469,HA_out_469}=HA_cout_391+HA_out_392;
  assign {HA_cout_470,HA_out_470}=HA_cout_392+HA_out_393;
  assign {HA_cout_471,HA_out_471}=HA_cout_393+HA_out_394;
  assign {HA_cout_472,HA_out_472}=HA_cout_394+HA_out_395;
  assign {HA_cout_473,HA_out_473}=HA_cout_395+HA_out_396;
  assign {HA_cout_474,HA_out_474}=HA_cout_396+HA_out_397;
  assign {HA_cout_475,HA_out_475}=HA_cout_397+HA_out_398;
  assign {HA_cout_476,HA_out_476}=HA_cout_398+HA_out_399;
  assign {HA_cout_477,HA_out_477}=HA_cout_399+FA_out_3800;
  assign {HA_cout_478,HA_out_478}=FA_cout_3800+FA_out_3801;
  assign {HA_cout_479,HA_out_479}=FA_cout_3801+FA_out_3802;
  assign {HA_cout_480,HA_out_480}=FA_cout_3802+FA_out_3803;
  assign {HA_cout_481,HA_out_481}=FA_cout_3803+FA_out_3804;
  assign {HA_cout_482,HA_out_482}=FA_cout_3804+FA_out_3805;
  assign {HA_cout_483,HA_out_483}=FA_cout_3805+FA_out_3806;
  assign {HA_cout_484,HA_out_484}=FA_cout_3806+FA_out_3807;
  assign {HA_cout_485,HA_out_485}=FA_cout_3807+FA_out_3808;
  assign {HA_cout_486,HA_out_486}=FA_cout_3808+FA_out_3809;
  assign {HA_cout_487,HA_out_487}=FA_cout_3809+FA_out_3810;
  assign {HA_cout_488,HA_out_488}=FA_cout_3810+FA_out_3811;
  assign {HA_cout_489,HA_out_489}=FA_cout_3811+FA_out_3812;
  assign {HA_cout_490,HA_out_490}=FA_cout_3812+FA_out_3813;
  assign {HA_cout_491,HA_out_491}=FA_cout_3813+FA_out_3814;
  assign {HA_cout_492,HA_out_492}=FA_cout_3814+FA_out_3815;
  assign {HA_cout_493,HA_out_493}=FA_cout_3815+FA_out_3816;
  assign {HA_cout_494,HA_out_494}=FA_cout_3816+FA_out_3817;
  assign {HA_cout_495,HA_out_495}=FA_cout_3817+FA_out_3818;
  assign {HA_cout_496,HA_out_496}=FA_cout_3818+FA_out_3819;
  assign {HA_cout_497,HA_out_497}=FA_cout_3819+FA_out_3820;
  assign {HA_cout_498,HA_out_498}=FA_cout_3821+FA_out_3822;
  assign {HA_cout_499,HA_out_499}=FA_cout_3822+FA_out_3823;
  assign {HA_cout_500,HA_out_500}=FA_cout_3823+FA_out_3824;
  assign {HA_cout_501,HA_out_501}=FA_cout_3824+FA_out_3825;
  assign {HA_cout_502,HA_out_502}=FA_cout_3825+FA_out_3826;
  assign {HA_cout_503,HA_out_503}=FA_cout_3826+FA_out_3827;
  assign {HA_cout_504,HA_out_504}=FA_cout_3827+FA_out_3828;
  assign {HA_cout_505,HA_out_505}=FA_cout_3828+FA_out_3829;
  assign {HA_cout_506,HA_out_506}=FA_cout_3829+FA_out_3830;
  assign {HA_cout_507,HA_out_507}=FA_cout_3830+FA_out_3831;
  assign {HA_cout_508,HA_out_508}=FA_cout_3831+FA_out_3832;
  assign {HA_cout_509,HA_out_509}=FA_cout_3832+FA_out_3833;
  assign {HA_cout_510,HA_out_510}=FA_cout_3833+FA_out_3834;
  assign {HA_cout_511,HA_out_511}=FA_cout_3834+FA_out_3835;
  assign {HA_cout_512,HA_out_512}=FA_cout_3835+FA_out_3836;
  assign {HA_cout_513,HA_out_513}=FA_cout_3836+FA_out_3837;
  assign {HA_cout_514,HA_out_514}=FA_cout_3837+FA_out_3838;
  assign {HA_cout_515,HA_out_515}=FA_cout_3838+FA_out_3839;
  assign {HA_cout_516,HA_out_516}=FA_cout_3839+FA_out_3840;
  assign {HA_cout_517,HA_out_517}=FA_cout_3840+FA_out_3841;
  assign {HA_cout_518,HA_out_518}=FA_cout_3841+FA_out_3842;
  assign {HA_cout_519,HA_out_519}=FA_cout_3842+HA_out_400;
  assign {HA_cout_520,HA_out_520}=HA_cout_400+HA_out_401;
  assign {HA_cout_521,HA_out_521}=HA_cout_401+HA_out_402;
  assign {HA_cout_522,HA_out_522}=HA_cout_402+HA_out_403;
  assign {HA_cout_523,HA_out_523}=HA_cout_403+HA_out_404;
  assign {HA_cout_524,HA_out_524}=HA_cout_404+HA_out_405;
  assign {HA_cout_525,HA_out_525}=HA_cout_405+HA_out_406;
  assign {HA_cout_526,HA_out_526}=HA_cout_406+HA_out_407;
  assign {HA_cout_527,HA_out_527}=HA_cout_407+HA_out_408;
  assign {HA_cout_528,HA_out_528}=HA_cout_408+HA_out_409;
  assign {HA_cout_529,HA_out_529}=HA_cout_409+HA_out_410;
  assign {HA_cout_530,HA_out_530}=HA_cout_410+HA_out_411;
  assign {HA_cout_531,HA_out_531}=HA_cout_411+HA_out_412;
  assign {HA_cout_532,HA_out_532}=HA_cout_412+HA_out_413;
  assign {HA_cout_533,HA_out_533}=HA_cout_413+HA_out_414;
  assign {HA_cout_534,HA_out_534}=HA_cout_414+HA_out_415;
  assign {HA_cout_535,HA_out_535}=HA_cout_415+HA_out_416;
  assign {HA_cout_536,HA_out_536}=HA_cout_416+HA_out_417;
  assign {HA_cout_537,HA_out_537}=HA_cout_417+HA_out_418;
  assign {HA_cout_538,HA_out_538}=HA_cout_418+HA_out_419;
  assign {HA_cout_539,HA_out_539}=HA_cout_419+HA_out_420;
  assign {HA_cout_540,HA_out_540}=HA_cout_420+HA_out_421;
  assign {HA_cout_541,HA_out_541}=HA_cout_421+HA_out_422;
  assign {HA_cout_542,HA_out_542}=HA_cout_422+HA_out_423;
  assign {HA_cout_543,HA_out_543}=HA_cout_423+HA_out_424;
  assign {HA_cout_544,HA_out_544}=HA_cout_424+HA_out_425;
  assign {HA_cout_545,HA_out_545}=HA_cout_425+HA_out_426;
  assign {HA_cout_546,HA_out_546}=HA_cout_426+HA_out_427;
  assign {HA_cout_547,HA_out_547}=HA_cout_427+HA_out_428;
  assign {HA_cout_548,HA_out_548}=HA_cout_428+HA_out_429;
  assign {HA_cout_549,HA_out_549}=HA_cout_429+HA_out_430;
  assign {HA_cout_550,HA_out_550}=HA_cout_430+HA_out_431;
  assign {HA_cout_551,HA_out_551}=HA_cout_431+HA_out_432;
  assign {HA_cout_552,HA_out_552}=HA_cout_432+HA_out_433;
  assign {HA_cout_553,HA_out_553}=HA_cout_433+HA_out_434;
  assign {HA_cout_554,HA_out_554}=HA_cout_434+HA_out_435;
  assign {HA_cout_555,HA_out_555}=HA_cout_435+HA_out_436;
  assign {HA_cout_556,HA_out_556}=HA_cout_436+HA_out_437;
  assign {HA_cout_557,HA_out_557}=HA_cout_437+HA_out_438;
  assign {HA_cout_558,HA_out_558}=HA_cout_438+HA_out_439;
  assign {HA_cout_559,HA_out_559}=HA_cout_439+HA_out_440;
  assign {HA_cout_560,HA_out_560}=HA_cout_440+REGS_1599;


  always @(negedge clk)
  begin
      REGS_0<=inp_0[0];
      REGS_1<=HA_out_0;
      REGS_2<=HA_out_42;
      REGS_3<=HA_out_84;
      REGS_4<=HA_cout_84;
      REGS_5<=HA_cout_85;
      REGS_6<=FA_cout_2205;
      REGS_7<=FA_cout_2206;
      REGS_8<=FA_cout_2207;
      REGS_9<=FA_cout_2208;
      REGS_10<=FA_cout_2209;
      REGS_11<=FA_cout_2210;
      REGS_12<=FA_cout_2211;
      REGS_13<=FA_cout_2212;
      REGS_14<=FA_cout_2213;
      REGS_15<=FA_cout_2214;
      REGS_16<=FA_cout_2215;
      REGS_17<=FA_cout_2216;
      REGS_18<=FA_cout_2217;
      REGS_19<=FA_cout_2218;
      REGS_20<=FA_cout_2219;
      REGS_21<=FA_cout_2220;
      REGS_22<=FA_cout_2221;
      REGS_23<=FA_cout_2222;
      REGS_24<=FA_cout_2223;
      REGS_25<=FA_cout_2224;
      REGS_26<=FA_cout_2225;
      REGS_27<=FA_cout_2226;
      REGS_28<=FA_cout_2227;
      REGS_29<=FA_cout_2228;
      REGS_30<=FA_cout_2229;
      REGS_31<=FA_cout_2230;
      REGS_32<=FA_cout_2231;
      REGS_33<=FA_cout_2232;
      REGS_34<=FA_cout_2233;
      REGS_35<=FA_cout_2234;
      REGS_36<=FA_cout_2235;
      REGS_37<=FA_cout_2236;
      REGS_38<=FA_cout_2237;
      REGS_39<=FA_cout_2238;
      REGS_40<=FA_cout_2239;
      REGS_41<=FA_cout_2240;
      REGS_42<=FA_cout_2241;
      REGS_43<=FA_cout_2242;
      REGS_44<=FA_cout_2243;
      REGS_45<=FA_cout_2244;
      REGS_46<=FA_cout_2245;
      REGS_47<=FA_cout_2246;
      REGS_48<=FA_cout_2247;
      REGS_49<=FA_cout_2248;
      REGS_50<=FA_cout_2249;
      REGS_51<=FA_cout_2250;
      REGS_52<=FA_cout_2251;
      REGS_53<=FA_cout_2252;
      REGS_54<=FA_cout_2253;
      REGS_55<=FA_cout_2254;
      REGS_56<=FA_cout_2255;
      REGS_57<=FA_cout_2256;
      REGS_58<=FA_cout_2257;
      REGS_59<=FA_cout_2258;
      REGS_60<=FA_cout_2259;
      REGS_61<=FA_cout_2260;
      REGS_62<=FA_cout_2261;
      REGS_63<=FA_cout_2262;
      REGS_64<=FA_cout_2263;
      REGS_65<=FA_cout_2264;
      REGS_66<=FA_cout_2265;
      REGS_67<=HA_out_85;
      REGS_68<=FA_out_2205;
      REGS_69<=FA_out_2206;
      REGS_70<=FA_out_2207;
      REGS_71<=FA_out_2208;
      REGS_72<=FA_out_2209;
      REGS_73<=FA_out_2210;
      REGS_74<=FA_out_2211;
      REGS_75<=FA_out_2212;
      REGS_76<=FA_out_2213;
      REGS_77<=FA_out_2214;
      REGS_78<=FA_out_2215;
      REGS_79<=FA_out_2216;
      REGS_80<=FA_out_2217;
      REGS_81<=FA_out_2218;
      REGS_82<=FA_out_2219;
      REGS_83<=FA_out_2220;
      REGS_84<=FA_out_2221;
      REGS_85<=FA_out_2222;
      REGS_86<=FA_out_2223;
      REGS_87<=FA_out_2224;
      REGS_88<=FA_out_2225;
      REGS_89<=FA_out_2226;
      REGS_90<=FA_out_2227;
      REGS_91<=FA_out_2228;
      REGS_92<=FA_out_2229;
      REGS_93<=FA_out_2230;
      REGS_94<=FA_out_2231;
      REGS_95<=FA_out_2232;
      REGS_96<=FA_out_2233;
      REGS_97<=FA_out_2234;
      REGS_98<=FA_out_2235;
      REGS_99<=FA_out_2236;
      REGS_100<=FA_out_2237;
      REGS_101<=FA_out_2238;
      REGS_102<=FA_out_2239;
      REGS_103<=FA_out_2240;
      REGS_104<=FA_out_2241;
      REGS_105<=FA_out_2242;
      REGS_106<=FA_out_2243;
      REGS_107<=FA_out_2244;
      REGS_108<=FA_out_2245;
      REGS_109<=FA_out_2246;
      REGS_110<=FA_out_2247;
      REGS_111<=FA_out_2248;
      REGS_112<=FA_out_2249;
      REGS_113<=FA_out_2250;
      REGS_114<=FA_out_2251;
      REGS_115<=FA_out_2252;
      REGS_116<=FA_out_2253;
      REGS_117<=FA_out_2254;
      REGS_118<=FA_out_2255;
      REGS_119<=FA_out_2256;
      REGS_120<=FA_out_2257;
      REGS_121<=FA_out_2258;
      REGS_122<=FA_out_2259;
      REGS_123<=FA_out_2260;
      REGS_124<=FA_out_2261;
      REGS_125<=FA_out_2262;
      REGS_126<=FA_out_2263;
      REGS_127<=FA_out_2264;
      REGS_128<=FA_out_2265;
      REGS_129<=FA_out_2266;
      REGS_130<=FA_cout_2266;
      REGS_131<=FA_out_2267;
      REGS_132<=FA_cout_2267;
      REGS_133<=FA_out_2268;
      REGS_134<=FA_cout_2268;
      REGS_135<=FA_out_2269;
      REGS_136<=FA_cout_2269;
      REGS_137<=HA_out_44;
      REGS_138<=FA_out_1388;
      REGS_139<=HA_out_86;
      REGS_140<=HA_cout_86;
      REGS_141<=HA_cout_87;
      REGS_142<=HA_cout_88;
      REGS_143<=FA_cout_2270;
      REGS_144<=FA_cout_2271;
      REGS_145<=FA_cout_2272;
      REGS_146<=FA_cout_2273;
      REGS_147<=FA_cout_2274;
      REGS_148<=FA_cout_2275;
      REGS_149<=FA_cout_2276;
      REGS_150<=FA_cout_2277;
      REGS_151<=FA_cout_2278;
      REGS_152<=FA_cout_2279;
      REGS_153<=FA_cout_2280;
      REGS_154<=FA_cout_2281;
      REGS_155<=FA_cout_2282;
      REGS_156<=FA_cout_2283;
      REGS_157<=FA_cout_2284;
      REGS_158<=FA_cout_2285;
      REGS_159<=FA_cout_2286;
      REGS_160<=FA_cout_2287;
      REGS_161<=FA_cout_2288;
      REGS_162<=FA_cout_2289;
      REGS_163<=FA_cout_2290;
      REGS_164<=FA_cout_2291;
      REGS_165<=FA_cout_2292;
      REGS_166<=FA_cout_2293;
      REGS_167<=FA_cout_2294;
      REGS_168<=FA_cout_2295;
      REGS_169<=FA_cout_2296;
      REGS_170<=FA_cout_2297;
      REGS_171<=FA_cout_2298;
      REGS_172<=FA_cout_2299;
      REGS_173<=FA_cout_2300;
      REGS_174<=FA_cout_2301;
      REGS_175<=FA_cout_2302;
      REGS_176<=FA_cout_2303;
      REGS_177<=FA_cout_2304;
      REGS_178<=FA_cout_2305;
      REGS_179<=FA_cout_2306;
      REGS_180<=FA_cout_2307;
      REGS_181<=FA_cout_2308;
      REGS_182<=FA_cout_2309;
      REGS_183<=FA_cout_2310;
      REGS_184<=FA_cout_2311;
      REGS_185<=FA_cout_2312;
      REGS_186<=FA_cout_2313;
      REGS_187<=FA_cout_2314;
      REGS_188<=FA_cout_2315;
      REGS_189<=FA_cout_2316;
      REGS_190<=FA_cout_2317;
      REGS_191<=FA_cout_2318;
      REGS_192<=FA_cout_2319;
      REGS_193<=FA_cout_2320;
      REGS_194<=FA_cout_2321;
      REGS_195<=FA_cout_2322;
      REGS_196<=FA_cout_2323;
      REGS_197<=FA_out_2324;
      REGS_198<=FA_cout_2324;
      REGS_199<=HA_out_87;
      REGS_200<=HA_out_88;
      REGS_201<=FA_out_2270;
      REGS_202<=FA_out_2271;
      REGS_203<=FA_out_2272;
      REGS_204<=FA_out_2273;
      REGS_205<=FA_out_2274;
      REGS_206<=FA_out_2275;
      REGS_207<=FA_out_2276;
      REGS_208<=FA_out_2277;
      REGS_209<=FA_out_2278;
      REGS_210<=FA_out_2279;
      REGS_211<=FA_out_2280;
      REGS_212<=FA_out_2281;
      REGS_213<=FA_out_2282;
      REGS_214<=FA_out_2283;
      REGS_215<=FA_out_2284;
      REGS_216<=FA_out_2285;
      REGS_217<=FA_out_2286;
      REGS_218<=FA_out_2287;
      REGS_219<=FA_out_2288;
      REGS_220<=FA_out_2289;
      REGS_221<=FA_out_2290;
      REGS_222<=FA_out_2291;
      REGS_223<=FA_out_2292;
      REGS_224<=FA_out_2293;
      REGS_225<=FA_out_2294;
      REGS_226<=FA_out_2295;
      REGS_227<=FA_out_2296;
      REGS_228<=FA_out_2297;
      REGS_229<=FA_out_2298;
      REGS_230<=FA_out_2299;
      REGS_231<=FA_out_2300;
      REGS_232<=FA_out_2301;
      REGS_233<=FA_out_2302;
      REGS_234<=FA_out_2303;
      REGS_235<=FA_out_2304;
      REGS_236<=FA_out_2305;
      REGS_237<=FA_out_2306;
      REGS_238<=FA_out_2307;
      REGS_239<=FA_out_2308;
      REGS_240<=FA_out_2309;
      REGS_241<=FA_out_2310;
      REGS_242<=FA_out_2311;
      REGS_243<=FA_out_2312;
      REGS_244<=FA_out_2313;
      REGS_245<=FA_out_2314;
      REGS_246<=FA_out_2315;
      REGS_247<=FA_out_2316;
      REGS_248<=FA_out_2317;
      REGS_249<=FA_out_2318;
      REGS_250<=FA_out_2319;
      REGS_251<=FA_out_2320;
      REGS_252<=FA_out_2321;
      REGS_253<=FA_out_2322;
      REGS_254<=FA_out_2323;
      REGS_255<=FA_out_2325;
      REGS_256<=FA_cout_2325;
      REGS_257<=FA_out_2326;
      REGS_258<=FA_cout_2326;
      REGS_259<=FA_out_2327;
      REGS_260<=FA_cout_2327;
      REGS_261<=FA_out_2328;
      REGS_262<=FA_cout_2328;
      REGS_263<=FA_out_2329;
      REGS_264<=FA_cout_2329;
      REGS_265<=FA_out_2330;
      REGS_266<=FA_cout_2330;
      REGS_267<=FA_out_2331;
      REGS_268<=FA_cout_2331;
      REGS_269<=FA_out_2332;
      REGS_270<=FA_cout_2332;
      REGS_271<=FA_out_2333;
      REGS_272<=FA_cout_2333;
      REGS_273<=FA_out_2334;
      REGS_274<=FA_cout_2334;
      REGS_275<=FA_out_2335;
      REGS_276<=FA_cout_2335;
      REGS_277<=FA_out_2336;
      REGS_278<=FA_cout_2336;
      REGS_279<=FA_out_2337;
      REGS_280<=FA_cout_2337;
      REGS_281<=FA_out_2338;
      REGS_282<=FA_cout_2338;
      REGS_283<=FA_out_256;
      REGS_284<=HA_out_46;
      REGS_285<=HA_out_89;
      REGS_286<=HA_cout_89;
      REGS_287<=HA_cout_90;
      REGS_288<=FA_cout_2339;
      REGS_289<=FA_cout_2340;
      REGS_290<=FA_cout_2341;
      REGS_291<=FA_cout_2342;
      REGS_292<=FA_cout_2343;
      REGS_293<=FA_cout_2344;
      REGS_294<=FA_cout_2345;
      REGS_295<=FA_cout_2346;
      REGS_296<=FA_cout_2347;
      REGS_297<=FA_cout_2348;
      REGS_298<=FA_cout_2349;
      REGS_299<=FA_cout_2350;
      REGS_300<=FA_cout_2351;
      REGS_301<=FA_cout_2352;
      REGS_302<=FA_cout_2353;
      REGS_303<=FA_cout_2354;
      REGS_304<=FA_cout_2355;
      REGS_305<=FA_cout_2356;
      REGS_306<=FA_cout_2357;
      REGS_307<=FA_cout_2358;
      REGS_308<=FA_cout_2359;
      REGS_309<=FA_cout_2360;
      REGS_310<=FA_cout_2361;
      REGS_311<=FA_cout_2362;
      REGS_312<=FA_cout_2363;
      REGS_313<=FA_cout_2364;
      REGS_314<=FA_cout_2365;
      REGS_315<=FA_cout_2366;
      REGS_316<=FA_cout_2367;
      REGS_317<=FA_cout_2368;
      REGS_318<=FA_cout_2369;
      REGS_319<=FA_cout_2370;
      REGS_320<=FA_cout_2371;
      REGS_321<=FA_cout_2372;
      REGS_322<=FA_cout_2373;
      REGS_323<=FA_cout_2374;
      REGS_324<=FA_cout_2375;
      REGS_325<=FA_cout_2376;
      REGS_326<=FA_cout_2377;
      REGS_327<=FA_cout_2378;
      REGS_328<=FA_cout_2379;
      REGS_329<=FA_cout_2380;
      REGS_330<=FA_cout_2381;
      REGS_331<=FA_cout_2382;
      REGS_332<=FA_cout_2383;
      REGS_333<=FA_cout_2384;
      REGS_334<=FA_cout_2385;
      REGS_335<=FA_cout_2386;
      REGS_336<=FA_out_2387;
      REGS_337<=FA_cout_2387;
      REGS_338<=FA_out_2388;
      REGS_339<=FA_cout_2388;
      REGS_340<=HA_out_90;
      REGS_341<=FA_out_2339;
      REGS_342<=FA_out_2340;
      REGS_343<=FA_out_2341;
      REGS_344<=FA_out_2342;
      REGS_345<=FA_out_2343;
      REGS_346<=FA_out_2344;
      REGS_347<=FA_out_2345;
      REGS_348<=FA_out_2346;
      REGS_349<=FA_out_2347;
      REGS_350<=FA_out_2348;
      REGS_351<=FA_out_2349;
      REGS_352<=FA_out_2350;
      REGS_353<=FA_out_2351;
      REGS_354<=FA_out_2352;
      REGS_355<=FA_out_2353;
      REGS_356<=FA_out_2354;
      REGS_357<=FA_out_2355;
      REGS_358<=FA_out_2356;
      REGS_359<=FA_out_2357;
      REGS_360<=FA_out_2358;
      REGS_361<=FA_out_2359;
      REGS_362<=FA_out_2360;
      REGS_363<=FA_out_2361;
      REGS_364<=FA_out_2362;
      REGS_365<=FA_out_2363;
      REGS_366<=FA_out_2364;
      REGS_367<=FA_out_2365;
      REGS_368<=FA_out_2366;
      REGS_369<=FA_out_2367;
      REGS_370<=FA_out_2368;
      REGS_371<=FA_out_2369;
      REGS_372<=FA_out_2370;
      REGS_373<=FA_out_2371;
      REGS_374<=FA_out_2372;
      REGS_375<=FA_out_2373;
      REGS_376<=FA_out_2374;
      REGS_377<=FA_out_2375;
      REGS_378<=FA_out_2376;
      REGS_379<=FA_out_2377;
      REGS_380<=FA_out_2378;
      REGS_381<=FA_out_2379;
      REGS_382<=FA_out_2380;
      REGS_383<=FA_out_2381;
      REGS_384<=FA_out_2382;
      REGS_385<=FA_out_2383;
      REGS_386<=FA_out_2384;
      REGS_387<=FA_out_2385;
      REGS_388<=FA_out_2386;
      REGS_389<=FA_out_2389;
      REGS_390<=FA_cout_2389;
      REGS_391<=FA_out_2390;
      REGS_392<=FA_cout_2390;
      REGS_393<=FA_out_2391;
      REGS_394<=FA_cout_2391;
      REGS_395<=FA_out_2392;
      REGS_396<=FA_cout_2392;
      REGS_397<=FA_out_2393;
      REGS_398<=FA_cout_2393;
      REGS_399<=FA_out_2394;
      REGS_400<=FA_cout_2394;
      REGS_401<=FA_out_2395;
      REGS_402<=FA_cout_2395;
      REGS_403<=FA_out_2396;
      REGS_404<=FA_cout_2396;
      REGS_405<=FA_out_2397;
      REGS_406<=FA_cout_2397;
      REGS_407<=FA_out_2398;
      REGS_408<=FA_cout_2398;
      REGS_409<=FA_out_2399;
      REGS_410<=FA_cout_2399;
      REGS_411<=FA_out_2400;
      REGS_412<=FA_cout_2400;
      REGS_413<=FA_out_2401;
      REGS_414<=FA_cout_2401;
      REGS_415<=FA_out_2402;
      REGS_416<=FA_cout_2402;
      REGS_417<=FA_out_2403;
      REGS_418<=FA_cout_2403;
      REGS_419<=FA_out_1585;
      REGS_420<=FA_out_1586;
      REGS_421<=HA_out_91;
      REGS_422<=HA_cout_91;
      REGS_423<=HA_cout_92;
      REGS_424<=FA_cout_2404;
      REGS_425<=FA_cout_2405;
      REGS_426<=FA_cout_2406;
      REGS_427<=FA_cout_2407;
      REGS_428<=FA_cout_2408;
      REGS_429<=FA_cout_2409;
      REGS_430<=FA_cout_2410;
      REGS_431<=FA_cout_2411;
      REGS_432<=FA_cout_2412;
      REGS_433<=FA_cout_2413;
      REGS_434<=FA_cout_2414;
      REGS_435<=FA_cout_2415;
      REGS_436<=FA_cout_2416;
      REGS_437<=FA_cout_2417;
      REGS_438<=FA_cout_2418;
      REGS_439<=FA_cout_2419;
      REGS_440<=FA_cout_2420;
      REGS_441<=FA_cout_2421;
      REGS_442<=FA_cout_2422;
      REGS_443<=FA_cout_2423;
      REGS_444<=FA_cout_2424;
      REGS_445<=FA_cout_2425;
      REGS_446<=FA_cout_2426;
      REGS_447<=FA_cout_2427;
      REGS_448<=FA_cout_2428;
      REGS_449<=FA_cout_2429;
      REGS_450<=FA_cout_2430;
      REGS_451<=FA_cout_2431;
      REGS_452<=FA_cout_2432;
      REGS_453<=FA_cout_2433;
      REGS_454<=FA_cout_2434;
      REGS_455<=FA_cout_2435;
      REGS_456<=FA_cout_2436;
      REGS_457<=FA_cout_2437;
      REGS_458<=FA_cout_2438;
      REGS_459<=FA_cout_2439;
      REGS_460<=FA_cout_2440;
      REGS_461<=FA_cout_2441;
      REGS_462<=FA_cout_2442;
      REGS_463<=FA_cout_2443;
      REGS_464<=FA_cout_2444;
      REGS_465<=FA_out_2445;
      REGS_466<=FA_cout_2445;
      REGS_467<=FA_out_2446;
      REGS_468<=FA_cout_2446;
      REGS_469<=FA_out_2447;
      REGS_470<=FA_cout_2447;
      REGS_471<=HA_out_92;
      REGS_472<=FA_out_2404;
      REGS_473<=FA_out_2405;
      REGS_474<=FA_out_2406;
      REGS_475<=FA_out_2407;
      REGS_476<=FA_out_2408;
      REGS_477<=FA_out_2409;
      REGS_478<=FA_out_2410;
      REGS_479<=FA_out_2411;
      REGS_480<=FA_out_2412;
      REGS_481<=FA_out_2413;
      REGS_482<=FA_out_2414;
      REGS_483<=FA_out_2415;
      REGS_484<=FA_out_2416;
      REGS_485<=FA_out_2417;
      REGS_486<=FA_out_2418;
      REGS_487<=FA_out_2419;
      REGS_488<=FA_out_2420;
      REGS_489<=FA_out_2421;
      REGS_490<=FA_out_2422;
      REGS_491<=FA_out_2423;
      REGS_492<=FA_out_2424;
      REGS_493<=FA_out_2425;
      REGS_494<=FA_out_2426;
      REGS_495<=FA_out_2427;
      REGS_496<=FA_out_2428;
      REGS_497<=FA_out_2429;
      REGS_498<=FA_out_2430;
      REGS_499<=FA_out_2431;
      REGS_500<=FA_out_2432;
      REGS_501<=FA_out_2433;
      REGS_502<=FA_out_2434;
      REGS_503<=FA_out_2435;
      REGS_504<=FA_out_2436;
      REGS_505<=FA_out_2437;
      REGS_506<=FA_out_2438;
      REGS_507<=FA_out_2439;
      REGS_508<=FA_out_2440;
      REGS_509<=FA_out_2441;
      REGS_510<=FA_out_2442;
      REGS_511<=FA_out_2443;
      REGS_512<=FA_out_2444;
      REGS_513<=FA_out_2448;
      REGS_514<=FA_cout_2448;
      REGS_515<=FA_out_2449;
      REGS_516<=FA_cout_2449;
      REGS_517<=FA_out_2450;
      REGS_518<=FA_cout_2450;
      REGS_519<=FA_out_2451;
      REGS_520<=FA_cout_2451;
      REGS_521<=FA_out_2452;
      REGS_522<=FA_cout_2452;
      REGS_523<=FA_out_2453;
      REGS_524<=FA_cout_2453;
      REGS_525<=FA_out_2454;
      REGS_526<=FA_cout_2454;
      REGS_527<=FA_out_2455;
      REGS_528<=FA_cout_2455;
      REGS_529<=FA_out_2456;
      REGS_530<=FA_cout_2456;
      REGS_531<=FA_out_2457;
      REGS_532<=FA_cout_2457;
      REGS_533<=FA_out_2458;
      REGS_534<=FA_cout_2458;
      REGS_535<=FA_out_2459;
      REGS_536<=FA_cout_2459;
      REGS_537<=FA_out_2460;
      REGS_538<=FA_cout_2460;
      REGS_539<=FA_out_2461;
      REGS_540<=FA_cout_2461;
      REGS_541<=FA_out_2462;
      REGS_542<=FA_cout_2462;
      REGS_543<=FA_out_2463;
      REGS_544<=FA_cout_2463;
      REGS_545<=FA_out_2464;
      REGS_546<=FA_cout_2464;
      REGS_547<=FA_out_2465;
      REGS_548<=FA_cout_2465;
      REGS_549<=FA_out_2466;
      REGS_550<=FA_cout_2466;
      REGS_551<=FA_out_2467;
      REGS_552<=FA_cout_2467;
      REGS_553<=FA_out_2468;
      REGS_554<=FA_cout_2468;
      REGS_555<=FA_out_2469;
      REGS_556<=FA_cout_2469;
      REGS_557<=FA_out_2470;
      REGS_558<=FA_cout_2470;
      REGS_559<=FA_out_2471;
      REGS_560<=FA_cout_2471;
      REGS_561<=FA_out_2472;
      REGS_562<=FA_cout_2472;
      REGS_563<=FA_out_2473;
      REGS_564<=FA_cout_2473;
      REGS_565<=FA_out_2474;
      REGS_566<=FA_cout_2474;
      REGS_567<=FA_out_2475;
      REGS_568<=FA_cout_2475;
      REGS_569<=inp_27[0];
      REGS_570<=HA_out_9;
      REGS_571<=HA_out_51;
      REGS_572<=HA_out_93;
      REGS_573<=HA_cout_93;
      REGS_574<=HA_cout_94;
      REGS_575<=FA_cout_2476;
      REGS_576<=FA_cout_2477;
      REGS_577<=FA_cout_2478;
      REGS_578<=FA_cout_2479;
      REGS_579<=FA_cout_2480;
      REGS_580<=FA_cout_2481;
      REGS_581<=FA_cout_2482;
      REGS_582<=FA_cout_2483;
      REGS_583<=FA_cout_2484;
      REGS_584<=FA_cout_2485;
      REGS_585<=FA_cout_2486;
      REGS_586<=FA_cout_2487;
      REGS_587<=FA_cout_2488;
      REGS_588<=FA_cout_2489;
      REGS_589<=FA_cout_2490;
      REGS_590<=FA_cout_2491;
      REGS_591<=FA_cout_2492;
      REGS_592<=FA_cout_2493;
      REGS_593<=FA_cout_2494;
      REGS_594<=FA_cout_2495;
      REGS_595<=FA_cout_2496;
      REGS_596<=FA_cout_2497;
      REGS_597<=FA_cout_2498;
      REGS_598<=FA_cout_2499;
      REGS_599<=FA_cout_2500;
      REGS_600<=FA_cout_2501;
      REGS_601<=FA_cout_2502;
      REGS_602<=FA_cout_2503;
      REGS_603<=FA_cout_2504;
      REGS_604<=FA_cout_2505;
      REGS_605<=FA_cout_2506;
      REGS_606<=FA_cout_2507;
      REGS_607<=FA_cout_2508;
      REGS_608<=FA_cout_2509;
      REGS_609<=FA_out_2510;
      REGS_610<=FA_cout_2510;
      REGS_611<=FA_out_2511;
      REGS_612<=FA_cout_2511;
      REGS_613<=FA_out_2512;
      REGS_614<=FA_cout_2512;
      REGS_615<=FA_out_2513;
      REGS_616<=FA_cout_2513;
      REGS_617<=HA_out_94;
      REGS_618<=FA_out_2476;
      REGS_619<=FA_out_2477;
      REGS_620<=FA_out_2478;
      REGS_621<=FA_out_2479;
      REGS_622<=FA_out_2480;
      REGS_623<=FA_out_2481;
      REGS_624<=FA_out_2482;
      REGS_625<=FA_out_2483;
      REGS_626<=FA_out_2484;
      REGS_627<=FA_out_2485;
      REGS_628<=FA_out_2486;
      REGS_629<=FA_out_2487;
      REGS_630<=FA_out_2488;
      REGS_631<=FA_out_2489;
      REGS_632<=FA_out_2490;
      REGS_633<=FA_out_2491;
      REGS_634<=FA_out_2492;
      REGS_635<=FA_out_2493;
      REGS_636<=FA_out_2494;
      REGS_637<=FA_out_2495;
      REGS_638<=FA_out_2496;
      REGS_639<=FA_out_2497;
      REGS_640<=FA_out_2498;
      REGS_641<=FA_out_2499;
      REGS_642<=FA_out_2500;
      REGS_643<=FA_out_2501;
      REGS_644<=FA_out_2502;
      REGS_645<=FA_out_2503;
      REGS_646<=FA_out_2504;
      REGS_647<=FA_out_2505;
      REGS_648<=FA_out_2506;
      REGS_649<=FA_out_2507;
      REGS_650<=FA_out_2508;
      REGS_651<=FA_out_2509;
      REGS_652<=FA_out_2514;
      REGS_653<=FA_cout_2514;
      REGS_654<=FA_out_2515;
      REGS_655<=FA_cout_2515;
      REGS_656<=FA_out_2516;
      REGS_657<=FA_cout_2516;
      REGS_658<=FA_out_2517;
      REGS_659<=FA_cout_2517;
      REGS_660<=FA_out_2518;
      REGS_661<=FA_cout_2518;
      REGS_662<=FA_out_2519;
      REGS_663<=FA_cout_2519;
      REGS_664<=FA_out_2520;
      REGS_665<=FA_cout_2520;
      REGS_666<=FA_out_2521;
      REGS_667<=FA_cout_2521;
      REGS_668<=FA_out_2522;
      REGS_669<=FA_cout_2522;
      REGS_670<=FA_out_2523;
      REGS_671<=FA_cout_2523;
      REGS_672<=FA_out_2524;
      REGS_673<=FA_cout_2524;
      REGS_674<=FA_out_2525;
      REGS_675<=FA_cout_2525;
      REGS_676<=FA_out_2526;
      REGS_677<=FA_cout_2526;
      REGS_678<=FA_out_2527;
      REGS_679<=FA_cout_2527;
      REGS_680<=FA_out_2528;
      REGS_681<=FA_cout_2528;
      REGS_682<=FA_out_2529;
      REGS_683<=FA_cout_2529;
      REGS_684<=FA_out_2530;
      REGS_685<=FA_cout_2530;
      REGS_686<=FA_out_2531;
      REGS_687<=FA_cout_2531;
      REGS_688<=FA_out_2532;
      REGS_689<=FA_cout_2532;
      REGS_690<=FA_out_2533;
      REGS_691<=FA_cout_2533;
      REGS_692<=HA_out_53;
      REGS_693<=FA_out_1778;
      REGS_694<=HA_out_95;
      REGS_695<=HA_cout_95;
      REGS_696<=HA_cout_96;
      REGS_697<=HA_cout_97;
      REGS_698<=FA_cout_2534;
      REGS_699<=FA_cout_2535;
      REGS_700<=FA_cout_2536;
      REGS_701<=FA_cout_2537;
      REGS_702<=FA_cout_2538;
      REGS_703<=FA_cout_2539;
      REGS_704<=FA_cout_2540;
      REGS_705<=FA_cout_2541;
      REGS_706<=FA_cout_2542;
      REGS_707<=FA_cout_2543;
      REGS_708<=FA_cout_2544;
      REGS_709<=FA_cout_2545;
      REGS_710<=FA_cout_2546;
      REGS_711<=FA_cout_2547;
      REGS_712<=FA_cout_2548;
      REGS_713<=FA_cout_2549;
      REGS_714<=FA_cout_2550;
      REGS_715<=FA_cout_2551;
      REGS_716<=FA_cout_2552;
      REGS_717<=FA_cout_2553;
      REGS_718<=FA_cout_2554;
      REGS_719<=FA_cout_2555;
      REGS_720<=FA_cout_2556;
      REGS_721<=FA_cout_2557;
      REGS_722<=FA_cout_2558;
      REGS_723<=FA_cout_2559;
      REGS_724<=FA_cout_2560;
      REGS_725<=FA_out_2561;
      REGS_726<=FA_cout_2561;
      REGS_727<=FA_out_2562;
      REGS_728<=FA_cout_2562;
      REGS_729<=FA_out_2563;
      REGS_730<=FA_cout_2563;
      REGS_731<=FA_out_2564;
      REGS_732<=FA_cout_2564;
      REGS_733<=FA_out_2565;
      REGS_734<=FA_cout_2565;
      REGS_735<=HA_out_96;
      REGS_736<=HA_out_97;
      REGS_737<=FA_out_2534;
      REGS_738<=FA_out_2535;
      REGS_739<=FA_out_2536;
      REGS_740<=FA_out_2537;
      REGS_741<=FA_out_2538;
      REGS_742<=FA_out_2539;
      REGS_743<=FA_out_2540;
      REGS_744<=FA_out_2541;
      REGS_745<=FA_out_2542;
      REGS_746<=FA_out_2543;
      REGS_747<=FA_out_2544;
      REGS_748<=FA_out_2545;
      REGS_749<=FA_out_2546;
      REGS_750<=FA_out_2547;
      REGS_751<=FA_out_2548;
      REGS_752<=FA_out_2549;
      REGS_753<=FA_out_2550;
      REGS_754<=FA_out_2551;
      REGS_755<=FA_out_2552;
      REGS_756<=FA_out_2553;
      REGS_757<=FA_out_2554;
      REGS_758<=FA_out_2555;
      REGS_759<=FA_out_2556;
      REGS_760<=FA_out_2557;
      REGS_761<=FA_out_2558;
      REGS_762<=FA_out_2559;
      REGS_763<=FA_out_2560;
      REGS_764<=FA_out_2566;
      REGS_765<=FA_cout_2566;
      REGS_766<=FA_out_2567;
      REGS_767<=FA_cout_2567;
      REGS_768<=FA_out_2568;
      REGS_769<=FA_cout_2568;
      REGS_770<=FA_out_2569;
      REGS_771<=FA_cout_2569;
      REGS_772<=FA_out_2570;
      REGS_773<=FA_cout_2570;
      REGS_774<=FA_out_2571;
      REGS_775<=FA_cout_2571;
      REGS_776<=FA_out_2572;
      REGS_777<=FA_cout_2572;
      REGS_778<=FA_out_2573;
      REGS_779<=FA_cout_2573;
      REGS_780<=FA_out_2574;
      REGS_781<=FA_cout_2574;
      REGS_782<=FA_out_2575;
      REGS_783<=FA_cout_2575;
      REGS_784<=FA_out_2576;
      REGS_785<=FA_cout_2576;
      REGS_786<=FA_out_2577;
      REGS_787<=FA_cout_2577;
      REGS_788<=FA_out_2578;
      REGS_789<=FA_cout_2578;
      REGS_790<=FA_out_2579;
      REGS_791<=FA_cout_2579;
      REGS_792<=FA_out_2580;
      REGS_793<=FA_cout_2580;
      REGS_794<=FA_out_2581;
      REGS_795<=FA_cout_2581;
      REGS_796<=FA_out_2582;
      REGS_797<=FA_cout_2582;
      REGS_798<=FA_out_2583;
      REGS_799<=FA_cout_2583;
      REGS_800<=FA_out_2584;
      REGS_801<=FA_cout_2584;
      REGS_802<=FA_out_2585;
      REGS_803<=FA_cout_2585;
      REGS_804<=FA_out_2586;
      REGS_805<=FA_cout_2586;
      REGS_806<=FA_out_2587;
      REGS_807<=FA_cout_2587;
      REGS_808<=FA_out_2588;
      REGS_809<=FA_cout_2588;
      REGS_810<=FA_out_2589;
      REGS_811<=FA_cout_2589;
      REGS_812<=FA_out_2590;
      REGS_813<=FA_cout_2590;
      REGS_814<=FA_out_2591;
      REGS_815<=FA_cout_2591;
      REGS_816<=FA_out_2592;
      REGS_817<=FA_cout_2592;
      REGS_818<=FA_out_2593;
      REGS_819<=FA_cout_2593;
      REGS_820<=FA_out_2594;
      REGS_821<=FA_cout_2594;
      REGS_822<=FA_out_2595;
      REGS_823<=FA_cout_2595;
      REGS_824<=FA_out_2596;
      REGS_825<=FA_cout_2596;
      REGS_826<=FA_out_2597;
      REGS_827<=FA_cout_2597;
      REGS_828<=FA_out_2598;
      REGS_829<=FA_cout_2598;
      REGS_830<=FA_out_2599;
      REGS_831<=FA_cout_2599;
      REGS_832<=FA_out_2600;
      REGS_833<=FA_cout_2600;
      REGS_834<=FA_out_2601;
      REGS_835<=FA_cout_2601;
      REGS_836<=FA_out_2602;
      REGS_837<=FA_cout_2602;
      REGS_838<=FA_out_2603;
      REGS_839<=FA_cout_2603;
      REGS_840<=FA_out_2604;
      REGS_841<=FA_cout_2604;
      REGS_842<=FA_out_2605;
      REGS_843<=FA_cout_2605;
      REGS_844<=FA_out_2606;
      REGS_845<=FA_cout_2606;
      REGS_846<=FA_out_2607;
      REGS_847<=FA_cout_2607;
      REGS_848<=FA_out_832;
      REGS_849<=HA_out_55;
      REGS_850<=HA_out_98;
      REGS_851<=HA_cout_98;
      REGS_852<=HA_cout_99;
      REGS_853<=FA_cout_2608;
      REGS_854<=FA_cout_2609;
      REGS_855<=FA_cout_2610;
      REGS_856<=FA_cout_2611;
      REGS_857<=FA_cout_2612;
      REGS_858<=FA_cout_2613;
      REGS_859<=FA_cout_2614;
      REGS_860<=FA_cout_2615;
      REGS_861<=FA_cout_2616;
      REGS_862<=FA_cout_2617;
      REGS_863<=FA_cout_2618;
      REGS_864<=FA_cout_2619;
      REGS_865<=FA_cout_2620;
      REGS_866<=FA_cout_2621;
      REGS_867<=FA_cout_2622;
      REGS_868<=FA_cout_2623;
      REGS_869<=FA_cout_2624;
      REGS_870<=FA_cout_2625;
      REGS_871<=FA_cout_2626;
      REGS_872<=FA_cout_2627;
      REGS_873<=FA_cout_2628;
      REGS_874<=FA_out_2629;
      REGS_875<=FA_cout_2629;
      REGS_876<=FA_out_2630;
      REGS_877<=FA_cout_2630;
      REGS_878<=FA_out_2631;
      REGS_879<=FA_cout_2631;
      REGS_880<=FA_out_2632;
      REGS_881<=FA_cout_2632;
      REGS_882<=FA_out_2633;
      REGS_883<=FA_cout_2633;
      REGS_884<=FA_out_2634;
      REGS_885<=FA_cout_2634;
      REGS_886<=HA_out_99;
      REGS_887<=FA_out_2608;
      REGS_888<=FA_out_2609;
      REGS_889<=FA_out_2610;
      REGS_890<=FA_out_2611;
      REGS_891<=FA_out_2612;
      REGS_892<=FA_out_2613;
      REGS_893<=FA_out_2614;
      REGS_894<=FA_out_2615;
      REGS_895<=FA_out_2616;
      REGS_896<=FA_out_2617;
      REGS_897<=FA_out_2618;
      REGS_898<=FA_out_2619;
      REGS_899<=FA_out_2620;
      REGS_900<=FA_out_2621;
      REGS_901<=FA_out_2622;
      REGS_902<=FA_out_2623;
      REGS_903<=FA_out_2624;
      REGS_904<=FA_out_2625;
      REGS_905<=FA_out_2626;
      REGS_906<=FA_out_2627;
      REGS_907<=FA_out_2628;
      REGS_908<=FA_out_2635;
      REGS_909<=FA_cout_2635;
      REGS_910<=FA_out_2636;
      REGS_911<=FA_cout_2636;
      REGS_912<=FA_out_2637;
      REGS_913<=FA_cout_2637;
      REGS_914<=FA_out_2638;
      REGS_915<=FA_cout_2638;
      REGS_916<=FA_out_2639;
      REGS_917<=FA_cout_2639;
      REGS_918<=FA_out_2640;
      REGS_919<=FA_cout_2640;
      REGS_920<=FA_out_2641;
      REGS_921<=FA_cout_2641;
      REGS_922<=FA_out_2642;
      REGS_923<=FA_cout_2642;
      REGS_924<=FA_out_2643;
      REGS_925<=FA_cout_2643;
      REGS_926<=FA_out_2644;
      REGS_927<=FA_cout_2644;
      REGS_928<=FA_out_2645;
      REGS_929<=FA_cout_2645;
      REGS_930<=FA_out_2646;
      REGS_931<=FA_cout_2646;
      REGS_932<=FA_out_2647;
      REGS_933<=FA_cout_2647;
      REGS_934<=FA_out_2648;
      REGS_935<=FA_cout_2648;
      REGS_936<=FA_out_2649;
      REGS_937<=FA_cout_2649;
      REGS_938<=FA_out_2650;
      REGS_939<=FA_cout_2650;
      REGS_940<=FA_out_2651;
      REGS_941<=FA_cout_2651;
      REGS_942<=FA_out_2652;
      REGS_943<=FA_cout_2652;
      REGS_944<=FA_out_2653;
      REGS_945<=FA_cout_2653;
      REGS_946<=FA_out_2654;
      REGS_947<=FA_cout_2654;
      REGS_948<=FA_out_2655;
      REGS_949<=FA_cout_2655;
      REGS_950<=FA_out_2656;
      REGS_951<=FA_cout_2656;
      REGS_952<=FA_out_2657;
      REGS_953<=FA_cout_2657;
      REGS_954<=FA_out_2658;
      REGS_955<=FA_cout_2658;
      REGS_956<=FA_out_2659;
      REGS_957<=FA_cout_2659;
      REGS_958<=FA_out_2660;
      REGS_959<=FA_cout_2660;
      REGS_960<=FA_out_2661;
      REGS_961<=FA_cout_2661;
      REGS_962<=FA_out_2662;
      REGS_963<=FA_cout_2662;
      REGS_964<=FA_out_2663;
      REGS_965<=FA_cout_2663;
      REGS_966<=FA_out_2664;
      REGS_967<=FA_cout_2664;
      REGS_968<=FA_out_2665;
      REGS_969<=FA_cout_2665;
      REGS_970<=FA_out_2666;
      REGS_971<=FA_cout_2666;
      REGS_972<=FA_out_2667;
      REGS_973<=FA_cout_2667;
      REGS_974<=FA_out_2668;
      REGS_975<=FA_cout_2668;
      REGS_976<=FA_out_2669;
      REGS_977<=FA_cout_2669;
      REGS_978<=FA_out_1978;
      REGS_979<=FA_out_1979;
      REGS_980<=HA_out_100;
      REGS_981<=HA_cout_100;
      REGS_982<=HA_cout_101;
      REGS_983<=FA_cout_2670;
      REGS_984<=FA_cout_2671;
      REGS_985<=FA_cout_2672;
      REGS_986<=FA_cout_2673;
      REGS_987<=FA_cout_2674;
      REGS_988<=FA_cout_2675;
      REGS_989<=FA_cout_2676;
      REGS_990<=FA_cout_2677;
      REGS_991<=FA_cout_2678;
      REGS_992<=FA_cout_2679;
      REGS_993<=FA_cout_2680;
      REGS_994<=FA_cout_2681;
      REGS_995<=FA_cout_2682;
      REGS_996<=FA_cout_2683;
      REGS_997<=FA_out_2684;
      REGS_998<=FA_cout_2684;
      REGS_999<=FA_out_2685;
      REGS_1000<=FA_cout_2685;
      REGS_1001<=FA_out_2686;
      REGS_1002<=FA_cout_2686;
      REGS_1003<=FA_out_2687;
      REGS_1004<=FA_cout_2687;
      REGS_1005<=FA_out_2688;
      REGS_1006<=FA_cout_2688;
      REGS_1007<=FA_out_2689;
      REGS_1008<=FA_cout_2689;
      REGS_1009<=FA_out_2690;
      REGS_1010<=FA_cout_2690;
      REGS_1011<=HA_out_101;
      REGS_1012<=FA_out_2670;
      REGS_1013<=FA_out_2671;
      REGS_1014<=FA_out_2672;
      REGS_1015<=FA_out_2673;
      REGS_1016<=FA_out_2674;
      REGS_1017<=FA_out_2675;
      REGS_1018<=FA_out_2676;
      REGS_1019<=FA_out_2677;
      REGS_1020<=FA_out_2678;
      REGS_1021<=FA_out_2679;
      REGS_1022<=FA_out_2680;
      REGS_1023<=FA_out_2681;
      REGS_1024<=FA_out_2682;
      REGS_1025<=FA_out_2683;
      REGS_1026<=FA_out_2691;
      REGS_1027<=FA_cout_2691;
      REGS_1028<=FA_out_2692;
      REGS_1029<=FA_cout_2692;
      REGS_1030<=FA_out_2693;
      REGS_1031<=FA_cout_2693;
      REGS_1032<=FA_out_2694;
      REGS_1033<=FA_cout_2694;
      REGS_1034<=FA_out_2695;
      REGS_1035<=FA_cout_2695;
      REGS_1036<=FA_out_2696;
      REGS_1037<=FA_cout_2696;
      REGS_1038<=FA_out_2697;
      REGS_1039<=FA_cout_2697;
      REGS_1040<=FA_out_2698;
      REGS_1041<=FA_cout_2698;
      REGS_1042<=FA_out_2699;
      REGS_1043<=FA_cout_2699;
      REGS_1044<=FA_out_2700;
      REGS_1045<=FA_cout_2700;
      REGS_1046<=FA_out_2701;
      REGS_1047<=FA_cout_2701;
      REGS_1048<=FA_out_2702;
      REGS_1049<=FA_cout_2702;
      REGS_1050<=FA_out_2703;
      REGS_1051<=FA_cout_2703;
      REGS_1052<=FA_out_2704;
      REGS_1053<=FA_cout_2704;
      REGS_1054<=FA_out_2705;
      REGS_1055<=FA_cout_2705;
      REGS_1056<=FA_out_2706;
      REGS_1057<=FA_cout_2706;
      REGS_1058<=FA_out_2707;
      REGS_1059<=FA_cout_2707;
      REGS_1060<=FA_out_2708;
      REGS_1061<=FA_cout_2708;
      REGS_1062<=FA_out_2709;
      REGS_1063<=FA_cout_2709;
      REGS_1064<=FA_out_2710;
      REGS_1065<=FA_cout_2710;
      REGS_1066<=FA_out_2711;
      REGS_1067<=FA_cout_2711;
      REGS_1068<=FA_out_2712;
      REGS_1069<=FA_cout_2712;
      REGS_1070<=FA_out_2713;
      REGS_1071<=FA_cout_2713;
      REGS_1072<=FA_out_2714;
      REGS_1073<=FA_cout_2714;
      REGS_1074<=FA_out_2715;
      REGS_1075<=FA_cout_2715;
      REGS_1076<=FA_out_2716;
      REGS_1077<=FA_cout_2716;
      REGS_1078<=FA_out_2717;
      REGS_1079<=FA_cout_2717;
      REGS_1080<=FA_out_2718;
      REGS_1081<=FA_cout_2718;
      REGS_1082<=FA_out_2719;
      REGS_1083<=FA_cout_2719;
      REGS_1084<=FA_out_2720;
      REGS_1085<=FA_cout_2720;
      REGS_1086<=FA_out_2721;
      REGS_1087<=FA_cout_2721;
      REGS_1088<=FA_out_2722;
      REGS_1089<=FA_cout_2722;
      REGS_1090<=FA_out_2723;
      REGS_1091<=FA_cout_2723;
      REGS_1092<=FA_out_2724;
      REGS_1093<=FA_cout_2724;
      REGS_1094<=FA_out_2725;
      REGS_1095<=FA_cout_2725;
      REGS_1096<=FA_out_2726;
      REGS_1097<=FA_cout_2726;
      REGS_1098<=FA_out_2727;
      REGS_1099<=FA_cout_2727;
      REGS_1100<=FA_out_2728;
      REGS_1101<=FA_cout_2728;
      REGS_1102<=FA_out_2729;
      REGS_1103<=FA_cout_2729;
      REGS_1104<=FA_out_2730;
      REGS_1105<=FA_cout_2730;
      REGS_1106<=FA_out_2731;
      REGS_1107<=FA_cout_2731;
      REGS_1108<=FA_out_2732;
      REGS_1109<=FA_cout_2732;
      REGS_1110<=FA_out_2733;
      REGS_1111<=FA_cout_2733;
      REGS_1112<=FA_out_2734;
      REGS_1113<=FA_cout_2734;
      REGS_1114<=FA_out_2735;
      REGS_1115<=FA_cout_2735;
      REGS_1116<=FA_out_2736;
      REGS_1117<=FA_cout_2736;
      REGS_1118<=FA_out_2737;
      REGS_1119<=FA_cout_2737;
      REGS_1120<=FA_out_2738;
      REGS_1121<=FA_cout_2738;
      REGS_1122<=FA_out_2739;
      REGS_1123<=FA_cout_2739;
      REGS_1124<=FA_out_2740;
      REGS_1125<=FA_cout_2740;
      REGS_1126<=FA_out_2741;
      REGS_1127<=FA_cout_2741;
      REGS_1128<=FA_out_2742;
      REGS_1129<=FA_cout_2742;
      REGS_1130<=FA_out_2743;
      REGS_1131<=FA_cout_2743;
      REGS_1132<=FA_out_2744;
      REGS_1133<=FA_cout_2744;
      REGS_1134<=FA_out_2745;
      REGS_1135<=FA_cout_2745;
      REGS_1136<=FA_out_2746;
      REGS_1137<=FA_cout_2746;
      REGS_1138<=inp_54[0];
      REGS_1139<=HA_out_18;
      REGS_1140<=HA_out_60;
      REGS_1141<=HA_out_102;
      REGS_1142<=HA_cout_102;
      REGS_1143<=HA_cout_103;
      REGS_1144<=FA_cout_2747;
      REGS_1145<=FA_cout_2748;
      REGS_1146<=FA_cout_2749;
      REGS_1147<=FA_cout_2750;
      REGS_1148<=FA_cout_2751;
      REGS_1149<=FA_cout_2752;
      REGS_1150<=FA_cout_2753;
      REGS_1151<=FA_out_2754;
      REGS_1152<=FA_cout_2754;
      REGS_1153<=FA_out_2755;
      REGS_1154<=FA_cout_2755;
      REGS_1155<=FA_out_2756;
      REGS_1156<=FA_cout_2756;
      REGS_1157<=FA_out_2757;
      REGS_1158<=FA_cout_2757;
      REGS_1159<=FA_out_2758;
      REGS_1160<=FA_cout_2758;
      REGS_1161<=FA_out_2759;
      REGS_1162<=FA_cout_2759;
      REGS_1163<=FA_out_2760;
      REGS_1164<=FA_cout_2760;
      REGS_1165<=FA_out_2761;
      REGS_1166<=FA_cout_2761;
      REGS_1167<=HA_out_103;
      REGS_1168<=FA_out_2747;
      REGS_1169<=FA_out_2748;
      REGS_1170<=FA_out_2749;
      REGS_1171<=FA_out_2750;
      REGS_1172<=FA_out_2751;
      REGS_1173<=FA_out_2752;
      REGS_1174<=FA_out_2753;
      REGS_1175<=FA_out_2762;
      REGS_1176<=FA_cout_2762;
      REGS_1177<=FA_out_2763;
      REGS_1178<=FA_cout_2763;
      REGS_1179<=FA_out_2764;
      REGS_1180<=FA_cout_2764;
      REGS_1181<=FA_out_2765;
      REGS_1182<=FA_cout_2765;
      REGS_1183<=FA_out_2766;
      REGS_1184<=FA_cout_2766;
      REGS_1185<=FA_out_2767;
      REGS_1186<=FA_cout_2767;
      REGS_1187<=FA_out_2768;
      REGS_1188<=FA_cout_2768;
      REGS_1189<=FA_out_2769;
      REGS_1190<=FA_cout_2769;
      REGS_1191<=FA_out_2770;
      REGS_1192<=FA_cout_2770;
      REGS_1193<=FA_out_2771;
      REGS_1194<=FA_cout_2771;
      REGS_1195<=FA_out_2772;
      REGS_1196<=FA_cout_2772;
      REGS_1197<=FA_out_2773;
      REGS_1198<=FA_cout_2773;
      REGS_1199<=FA_out_2774;
      REGS_1200<=FA_cout_2774;
      REGS_1201<=FA_out_2775;
      REGS_1202<=FA_cout_2775;
      REGS_1203<=FA_out_2776;
      REGS_1204<=FA_cout_2776;
      REGS_1205<=FA_out_2777;
      REGS_1206<=FA_cout_2777;
      REGS_1207<=FA_out_2778;
      REGS_1208<=FA_cout_2778;
      REGS_1209<=FA_out_2779;
      REGS_1210<=FA_cout_2779;
      REGS_1211<=FA_out_2780;
      REGS_1212<=FA_cout_2780;
      REGS_1213<=FA_out_2781;
      REGS_1214<=FA_cout_2781;
      REGS_1215<=FA_out_2782;
      REGS_1216<=FA_cout_2782;
      REGS_1217<=FA_out_2783;
      REGS_1218<=FA_cout_2783;
      REGS_1219<=FA_out_2784;
      REGS_1220<=FA_cout_2784;
      REGS_1221<=FA_out_2785;
      REGS_1222<=FA_cout_2785;
      REGS_1223<=FA_out_2786;
      REGS_1224<=FA_cout_2786;
      REGS_1225<=FA_out_2787;
      REGS_1226<=FA_cout_2787;
      REGS_1227<=FA_out_2788;
      REGS_1228<=FA_cout_2788;
      REGS_1229<=FA_out_2789;
      REGS_1230<=FA_cout_2789;
      REGS_1231<=HA_out_104;
      REGS_1232<=HA_cout_104;
      REGS_1233<=HA_out_105;
      REGS_1234<=HA_cout_105;
      REGS_1235<=HA_out_106;
      REGS_1236<=HA_cout_106;
      REGS_1237<=FA_out_2790;
      REGS_1238<=FA_cout_2790;
      REGS_1239<=HA_out_107;
      REGS_1240<=HA_cout_107;
      REGS_1241<=HA_out_108;
      REGS_1242<=HA_cout_108;
      REGS_1243<=HA_out_109;
      REGS_1244<=HA_cout_109;
      REGS_1245<=FA_out_2791;
      REGS_1246<=FA_cout_2791;
      REGS_1247<=HA_out_62;
      REGS_1248<=FA_out_2168;
      REGS_1249<=HA_out_110;
      REGS_1250<=HA_cout_110;
      REGS_1251<=FA_out_2184;
      REGS_1252<=HA_out_111;
      REGS_1253<=HA_cout_111;
      REGS_1254<=HA_out_112;
      REGS_1255<=HA_cout_112;
      REGS_1256<=HA_out_113;
      REGS_1257<=HA_cout_113;
      REGS_1258<=FA_out_2190;
      REGS_1259<=HA_out_114;
      REGS_1260<=HA_cout_114;
      REGS_1261<=HA_out_115;
      REGS_1262<=HA_cout_115;
      REGS_1263<=HA_out_116;
      REGS_1264<=HA_cout_116;
      REGS_1265<=FA_out_2196;
      REGS_1266<=HA_out_117;
      REGS_1267<=HA_cout_117;
      REGS_1268<=FA_out_2170;
      REGS_1269<=FA_out_2198;
      REGS_1270<=HA_out_118;
      REGS_1271<=HA_cout_118;
      REGS_1272<=HA_out_64;
      REGS_1273<=HA_out_119;
      REGS_1274<=HA_cout_119;
      REGS_1275<=FA_out_2201;
      REGS_1276<=HA_out_120;
      REGS_1277<=HA_cout_120;
      REGS_1278<=HA_out_67;
      REGS_1279<=HA_out_121;
      REGS_1280<=HA_cout_121;
      REGS_1281<=FA_out_2204;
      REGS_1282<=HA_out_122;
      REGS_1283<=HA_cout_122;
      REGS_1284<=FA_out_1303;
      REGS_1285<=HA_out_123;
      REGS_1286<=HA_cout_123;
      REGS_1287<=HA_out_71;
      REGS_1288<=FA_out_1312;
      REGS_1289<=HA_out_124;
      REGS_1290<=HA_cout_124;
      REGS_1291<=HA_out_74;
      REGS_1292<=FA_out_1321;
      REGS_1293<=HA_out_125;
      REGS_1294<=HA_cout_125;
      REGS_1295<=HA_cout_77;
      REGS_1296<=HA_out_78;
      REGS_1297<=HA_out_28;
      REGS_1298<=HA_cout_80;
      REGS_1299<=HA_out_81;
      REGS_1300<=HA_out_37;
      REGS_1301<=HA_cout_83;
      REGS_1302<=inp_63[24];
      REGS_1303<=inp_63[51];
      REGS_1304<=REGS_0;
      REGS_1305<=REGS_1;
      REGS_1306<=REGS_2;
      REGS_1307<=REGS_3;
      REGS_1308<=HA_out_126;
      REGS_1309<=HA_out_167;
      REGS_1310<=HA_out_209;
      REGS_1311<=HA_out_262;
      REGS_1312<=HA_out_310;
      REGS_1313<=HA_cout_310;
      REGS_1314<=HA_cout_311;
      REGS_1315<=HA_cout_312;
      REGS_1316<=HA_cout_313;
      REGS_1317<=HA_cout_314;
      REGS_1318<=HA_cout_315;
      REGS_1319<=HA_cout_316;
      REGS_1320<=HA_cout_317;
      REGS_1321<=HA_cout_318;
      REGS_1322<=HA_cout_319;
      REGS_1323<=HA_cout_320;
      REGS_1324<=HA_cout_321;
      REGS_1325<=HA_cout_322;
      REGS_1326<=HA_cout_323;
      REGS_1327<=HA_cout_324;
      REGS_1328<=HA_cout_325;
      REGS_1329<=HA_cout_326;
      REGS_1330<=HA_cout_327;
      REGS_1331<=HA_cout_328;
      REGS_1332<=HA_cout_329;
      REGS_1333<=HA_cout_330;
      REGS_1334<=HA_cout_331;
      REGS_1335<=HA_cout_332;
      REGS_1336<=HA_cout_333;
      REGS_1337<=FA_cout_3730;
      REGS_1338<=FA_cout_3731;
      REGS_1339<=FA_cout_3732;
      REGS_1340<=FA_cout_3733;
      REGS_1341<=FA_cout_3734;
      REGS_1342<=FA_cout_3735;
      REGS_1343<=FA_cout_3736;
      REGS_1344<=FA_cout_3737;
      REGS_1345<=FA_cout_3738;
      REGS_1346<=FA_cout_3739;
      REGS_1347<=FA_cout_3740;
      REGS_1348<=FA_cout_3741;
      REGS_1349<=FA_cout_3742;
      REGS_1350<=FA_cout_3743;
      REGS_1351<=FA_cout_3744;
      REGS_1352<=FA_cout_3745;
      REGS_1353<=FA_cout_3746;
      REGS_1354<=FA_cout_3747;
      REGS_1355<=FA_cout_3748;
      REGS_1356<=FA_cout_3749;
      REGS_1357<=FA_cout_3750;
      REGS_1358<=FA_cout_3751;
      REGS_1359<=FA_cout_3752;
      REGS_1360<=FA_cout_3753;
      REGS_1361<=FA_cout_3754;
      REGS_1362<=FA_cout_3755;
      REGS_1363<=FA_cout_3756;
      REGS_1364<=FA_cout_3757;
      REGS_1365<=FA_cout_3758;
      REGS_1366<=FA_cout_3759;
      REGS_1367<=FA_cout_3760;
      REGS_1368<=FA_cout_3761;
      REGS_1369<=FA_cout_3762;
      REGS_1370<=FA_cout_3763;
      REGS_1371<=FA_cout_3764;
      REGS_1372<=FA_cout_3765;
      REGS_1373<=FA_cout_3766;
      REGS_1374<=FA_cout_3767;
      REGS_1375<=FA_cout_3768;
      REGS_1376<=HA_out_311;
      REGS_1377<=HA_out_312;
      REGS_1378<=HA_out_313;
      REGS_1379<=HA_out_314;
      REGS_1380<=HA_out_315;
      REGS_1381<=HA_out_316;
      REGS_1382<=HA_out_317;
      REGS_1383<=HA_out_318;
      REGS_1384<=HA_out_319;
      REGS_1385<=HA_out_320;
      REGS_1386<=HA_out_321;
      REGS_1387<=HA_out_322;
      REGS_1388<=HA_out_323;
      REGS_1389<=HA_out_324;
      REGS_1390<=HA_out_325;
      REGS_1391<=HA_out_326;
      REGS_1392<=HA_out_327;
      REGS_1393<=HA_out_328;
      REGS_1394<=HA_out_329;
      REGS_1395<=HA_out_330;
      REGS_1396<=HA_out_331;
      REGS_1397<=HA_out_332;
      REGS_1398<=HA_out_333;
      REGS_1399<=FA_out_3730;
      REGS_1400<=FA_out_3731;
      REGS_1401<=FA_out_3732;
      REGS_1402<=FA_out_3733;
      REGS_1403<=FA_out_3734;
      REGS_1404<=FA_out_3735;
      REGS_1405<=FA_out_3736;
      REGS_1406<=FA_out_3737;
      REGS_1407<=FA_out_3738;
      REGS_1408<=FA_out_3739;
      REGS_1409<=FA_out_3740;
      REGS_1410<=FA_out_3741;
      REGS_1411<=FA_out_3742;
      REGS_1412<=FA_out_3743;
      REGS_1413<=FA_out_3744;
      REGS_1414<=FA_out_3745;
      REGS_1415<=FA_out_3746;
      REGS_1416<=FA_out_3747;
      REGS_1417<=FA_out_3748;
      REGS_1418<=FA_out_3749;
      REGS_1419<=FA_out_3750;
      REGS_1420<=FA_out_3751;
      REGS_1421<=FA_out_3752;
      REGS_1422<=FA_out_3753;
      REGS_1423<=FA_out_3754;
      REGS_1424<=FA_out_3755;
      REGS_1425<=FA_out_3756;
      REGS_1426<=FA_out_3757;
      REGS_1427<=FA_out_3758;
      REGS_1428<=FA_out_3759;
      REGS_1429<=FA_out_3760;
      REGS_1430<=FA_out_3761;
      REGS_1431<=FA_out_3762;
      REGS_1432<=FA_out_3763;
      REGS_1433<=FA_out_3764;
      REGS_1434<=FA_out_3765;
      REGS_1435<=FA_out_3766;
      REGS_1436<=FA_out_3767;
      REGS_1437<=FA_out_3768;
      REGS_1438<=FA_out_3769;
      REGS_1439<=FA_cout_3769;
      REGS_1440<=FA_out_3770;
      REGS_1441<=FA_cout_3770;
      REGS_1442<=FA_out_3771;
      REGS_1443<=FA_cout_3771;
      REGS_1444<=FA_out_3772;
      REGS_1445<=FA_cout_3772;
      REGS_1446<=FA_out_3773;
      REGS_1447<=FA_cout_3773;
      REGS_1448<=FA_out_3774;
      REGS_1449<=FA_cout_3774;
      REGS_1450<=FA_out_3775;
      REGS_1451<=FA_cout_3775;
      REGS_1452<=FA_out_3776;
      REGS_1453<=FA_cout_3776;
      REGS_1454<=FA_out_3777;
      REGS_1455<=FA_cout_3777;
      REGS_1456<=HA_out_278;
      REGS_1457<=HA_out_279;
      REGS_1458<=HA_out_280;
      REGS_1459<=HA_out_281;
      REGS_1460<=HA_out_282;
      REGS_1461<=HA_out_283;
      REGS_1462<=HA_out_284;
      REGS_1463<=FA_out_3669;
      REGS_1464<=FA_out_3670;
      REGS_1465<=FA_out_3671;
      REGS_1466<=FA_out_3672;
      REGS_1467<=FA_out_3673;
      REGS_1468<=FA_out_3674;
      REGS_1469<=FA_out_3675;
      REGS_1470<=FA_out_3676;
      REGS_1471<=FA_out_3677;
      REGS_1472<=FA_out_3678;
      REGS_1473<=FA_out_3679;
      REGS_1474<=FA_out_3680;
      REGS_1475<=FA_out_3681;
      REGS_1476<=HA_out_334;
      REGS_1477<=HA_cout_334;
      REGS_1478<=FA_out_3684;
      REGS_1479<=FA_out_3685;
      REGS_1480<=FA_out_3687;
      REGS_1481<=FA_out_3778;
      REGS_1482<=FA_cout_3778;
      REGS_1483<=FA_out_3683;
      REGS_1484<=FA_out_3689;
      REGS_1485<=FA_out_3779;
      REGS_1486<=FA_cout_3779;
      REGS_1487<=FA_out_3691;
      REGS_1488<=FA_out_3780;
      REGS_1489<=FA_cout_3780;
      REGS_1490<=FA_out_3693;
      REGS_1491<=FA_out_3781;
      REGS_1492<=FA_cout_3781;
      REGS_1493<=FA_out_3695;
      REGS_1494<=FA_out_3782;
      REGS_1495<=FA_cout_3782;
      REGS_1496<=FA_out_3697;
      REGS_1497<=FA_out_3783;
      REGS_1498<=FA_cout_3783;
      REGS_1499<=FA_out_3699;
      REGS_1500<=FA_out_3784;
      REGS_1501<=FA_cout_3784;
      REGS_1502<=FA_out_3701;
      REGS_1503<=FA_out_3785;
      REGS_1504<=FA_cout_3785;
      REGS_1505<=FA_out_3703;
      REGS_1506<=FA_out_3786;
      REGS_1507<=FA_cout_3786;
      REGS_1508<=FA_out_3705;
      REGS_1509<=FA_out_3787;
      REGS_1510<=FA_cout_3787;
      REGS_1511<=FA_out_3707;
      REGS_1512<=FA_out_3788;
      REGS_1513<=FA_cout_3788;
      REGS_1514<=FA_out_3709;
      REGS_1515<=FA_out_3789;
      REGS_1516<=FA_cout_3789;
      REGS_1517<=HA_out_285;
      REGS_1518<=FA_out_3790;
      REGS_1519<=FA_cout_3790;
      REGS_1520<=HA_out_286;
      REGS_1521<=FA_out_3791;
      REGS_1522<=FA_cout_3791;
      REGS_1523<=HA_out_287;
      REGS_1524<=FA_out_3792;
      REGS_1525<=FA_cout_3792;
      REGS_1526<=HA_out_288;
      REGS_1527<=FA_out_3793;
      REGS_1528<=FA_cout_3793;
      REGS_1529<=HA_out_289;
      REGS_1530<=FA_out_3794;
      REGS_1531<=FA_cout_3794;
      REGS_1532<=HA_out_290;
      REGS_1533<=FA_out_3795;
      REGS_1534<=FA_cout_3795;
      REGS_1535<=FA_out_3577;
      REGS_1536<=FA_out_3796;
      REGS_1537<=FA_cout_3796;
      REGS_1538<=FA_out_3797;
      REGS_1539<=FA_cout_3797;
      REGS_1540<=FA_out_3798;
      REGS_1541<=FA_cout_3798;
      REGS_1542<=FA_out_3799;
      REGS_1543<=FA_cout_3799;
      REGS_1544<=HA_out_335;
      REGS_1545<=HA_cout_335;
      REGS_1546<=HA_out_336;
      REGS_1547<=HA_cout_336;
      REGS_1548<=HA_out_337;
      REGS_1549<=HA_cout_337;
      REGS_1550<=HA_out_338;
      REGS_1551<=HA_cout_338;
      REGS_1552<=HA_out_339;
      REGS_1553<=HA_cout_339;
      REGS_1554<=HA_out_340;
      REGS_1555<=HA_cout_340;
      REGS_1556<=HA_out_341;
      REGS_1557<=HA_cout_341;
      REGS_1558<=HA_out_342;
      REGS_1559<=HA_cout_342;
      REGS_1560<=HA_out_343;
      REGS_1561<=HA_cout_343;
      REGS_1562<=HA_out_344;
      REGS_1563<=HA_cout_344;
      REGS_1564<=HA_out_345;
      REGS_1565<=HA_cout_345;
      REGS_1566<=HA_out_346;
      REGS_1567<=HA_cout_346;
      REGS_1568<=HA_out_347;
      REGS_1569<=HA_cout_347;
      REGS_1570<=HA_out_348;
      REGS_1571<=HA_cout_348;
      REGS_1572<=HA_out_349;
      REGS_1573<=HA_cout_349;
      REGS_1574<=HA_out_350;
      REGS_1575<=HA_cout_350;
      REGS_1576<=HA_out_351;
      REGS_1577<=HA_cout_351;
      REGS_1578<=HA_out_352;
      REGS_1579<=HA_cout_352;
      REGS_1580<=HA_out_353;
      REGS_1581<=HA_cout_353;
      REGS_1582<=HA_out_354;
      REGS_1583<=HA_cout_354;
      REGS_1584<=HA_out_355;
      REGS_1585<=HA_cout_355;
      REGS_1586<=HA_out_356;
      REGS_1587<=HA_cout_356;
      REGS_1588<=HA_out_357;
      REGS_1589<=HA_cout_357;
      REGS_1590<=HA_out_358;
      REGS_1591<=HA_cout_358;
      REGS_1592<=HA_out_359;
      REGS_1593<=HA_cout_359;
      REGS_1594<=HA_out_360;
      REGS_1595<=HA_cout_360;
      REGS_1596<=HA_out_361;
      REGS_1597<=HA_cout_361;
      REGS_1598<=HA_out_362;
      REGS_1599<=HA_cout_362;
  end


endmodule

