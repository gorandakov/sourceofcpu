/*
Copyright 2022-2024 Goran Dakov, see additional restriction in copying.txt

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/


`include "../struct.sv"

module normalizeD(
  clk,
  rst,
  A,
  isDBL,
  isEXT,
  en,
  clkEn,
  res
  );

  localparam [11:0] DEN_DBL=12'h400;
  localparam [15:0] DEN_EXT=16'h4000;
  input clk;
  input rst;
  input [81:0] A;
  input isDBL;
  input isEXT;
  input en;
  input clkEn;
  output [81:0] res;

  wire [15:0] expA;
  wire [15:0] denor_from;
  wire [15:0] offset;
  reg [15:0] offset_reg;

  assign expA=isDBL ? {A[65],{4{~A[65]}},A[63:53]} : {A[65],A[80:66]};
  assign denor_from=isDBL ? {DEN_DBL[11],{4{~DEN_DBL[11]}},DEN_DBL[10:0]} : DEN_EXT;

  adder #(16) offAdd_mod(denor_from,~expA,offset,1'b1,1'b1);

  generate
    genvar t;
    for(t=0;t<8;t=t+1) begin
	get_carry #(3) cmpUP_mod(offset_reg[5:3],~t[2:0],1'b1,coUP[t]);
	get_carry #(3) cmpDN_mod(offset_reg[2:0],~t[2:0],1'b1,coDN[t]);
	assign eqUP[t]=t==offset_reg[5:3];
	assign the_mask[8*t+:8]=~eqUP[t] & coUP[t] ? 8'b0 : 8'bz;
	assign the_mask[8*t+:8]=eqUP[t] ? submask : 8'bz;
	assign the_mask[8*t+:8]=~coUP[t] ? 8'hff : 8'bz
	assign submask[t]=coDN[t];
    end
  endgenerate
endmodule
