`define exc_gpf 0
`define exc_pf 1

