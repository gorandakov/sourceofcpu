operations.v