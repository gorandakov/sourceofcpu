/*
Copyright 2022 Goran Dakov

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

`include "struct.sv"


module DFF(clk,en,d,q);
  parameter WIDTH=1;
  input clk;
  input en;
  input [WIDTH-1:0] d;
  output reg [WIDTH-1:0] q;//={WIDTH{1'b0}};
  
  always @(posedge clk)
    begin
      if (en) q<=d;
    end

endmodule



module DFF2(clk,rst,en,d,q);
  parameter WIDTH=1;
  input clk;
  input rst;
  input en;
  input [WIDTH-1:0] d;
  output reg [WIDTH-1:0] q;//={WIDTH{1'b0}};
  
  always @(posedge clk)
    begin
	  if (rst) q<={WIDTH{1'B0}};
      else if (en) q<=d;
    end

endmodule


module muxx3(out,hitA,wf,inA,inB,inF);

  parameter WIDTH=1;

  output [WIDTH-1:0] out;
  input hitA;
  input wf;
  input [WIDTH-1:0] inA;
  input [WIDTH-1:0] inB;
  input [WIDTH-1:0] inF;

  assign out=(hitA & ~wf) ? inA : {WIDTH{{1{1'bz}}}};
  assign out=(~hitA & ~wf) ? inB : {WIDTH{{1{1'bz}}}};
  assign out=wf ? inF : {WIDTH{{1{1'bz}}}};

endmodule


module optional_register(
  clk,
  dataIn,dataOut);
  parameter WIDTH=32;
  parameter CNT=0;
  
  input clk;
  input  [WIDTH-1:0] dataIn;
  output [WIDTH-1:0] dataOut;
  
  reg [WIDTH-1:0] first;
  reg [WIDTH-1:0] second;

  always @(posedge clk) begin
      first<=dataIn;
      second<=first;
  end  

  generate
      if (CNT==0) assign dataOut=dataIn;
      if (CNT==1) assign dataOut=first;
      if (CNT==2) assign dataOut=second;
  endgenerate
  
endmodule

