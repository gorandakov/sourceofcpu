//comment for 128k cache
`define ICACHE_256K
//comment for 128k cache
`define DCACHE_256K
