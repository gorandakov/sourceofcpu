csrss_no.v