struct.v