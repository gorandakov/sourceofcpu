fpoperations.v